
module mult24_unsigned ( A, B, Z);
   input [23:0] A;
   input [23:0] B;
   output [47:0] Z;

   // Internal wires
   wire n_0;
   wire n_2;
   wire n_3;
   wire n_4;
   wire n_5;
   wire n_6;
   wire n_7;
   wire n_8;
   wire n_9;
   wire n_10;
   wire n_11;
   wire n_12;
   wire n_13;
   wire n_14;
   wire n_15;
   wire n_16;
   wire n_17;
   wire n_18;
   wire n_19;
   wire n_20;
   wire n_21;
   wire n_22;
   wire n_23;
   wire n_24;
   wire n_25;
   wire n_26;
   wire n_27;
   wire n_28;
   wire n_29;
   wire n_30;
   wire n_31;
   wire n_32;
   wire n_33;
   wire n_34;
   wire n_35;
   wire n_36;
   wire n_37;
   wire n_38;
   wire n_39;
   wire n_40;
   wire n_41;
   wire n_42;
   wire n_43;
   wire n_44;
   wire n_45;
   wire n_46;
   wire n_47;
   wire n_48;
   wire n_49;
   wire n_50;
   wire n_51;
   wire n_52;
   wire n_53;
   wire n_54;
   wire n_55;
   wire n_56;
   wire n_57;
   wire n_58;
   wire n_59;
   wire n_60;
   wire n_61;
   wire n_62;
   wire n_63;
   wire n_64;
   wire n_65;
   wire n_66;
   wire n_67;
   wire n_68;
   wire n_69;
   wire n_70;
   wire n_71;
   wire n_72;
   wire n_73;
   wire n_74;
   wire n_75;
   wire n_76;
   wire n_77;
   wire n_78;
   wire n_79;
   wire n_80;
   wire n_81;
   wire n_82;
   wire n_83;
   wire n_84;
   wire n_85;
   wire n_86;
   wire n_87;
   wire n_88;
   wire n_90;
   wire n_91;
   wire n_92;
   wire n_93;
   wire n_94;
   wire n_95;
   wire n_96;
   wire n_97;
   wire n_98;
   wire n_99;
   wire n_100;
   wire n_101;
   wire n_102;
   wire n_103;
   wire n_104;
   wire n_105;
   wire n_106;
   wire n_107;
   wire n_108;
   wire n_109;
   wire n_110;
   wire n_111;
   wire n_112;
   wire n_113;
   wire n_114;
   wire n_115;
   wire n_116;
   wire n_117;
   wire n_118;
   wire n_119;
   wire n_120;
   wire n_121;
   wire n_122;
   wire n_123;
   wire n_124;
   wire n_125;
   wire n_126;
   wire n_127;
   wire n_128;
   wire n_129;
   wire n_130;
   wire n_131;
   wire n_132;
   wire n_133;
   wire n_134;
   wire n_135;
   wire n_136;
   wire n_137;
   wire n_138;
   wire n_139;
   wire n_140;
   wire n_141;
   wire n_142;
   wire n_143;
   wire n_144;
   wire n_145;
   wire n_146;
   wire n_147;
   wire n_148;
   wire n_149;
   wire n_150;
   wire n_151;
   wire n_152;
   wire n_153;
   wire n_154;
   wire n_155;
   wire n_156;
   wire n_157;
   wire n_158;
   wire n_159;
   wire n_160;
   wire n_161;
   wire n_162;
   wire n_163;
   wire n_164;
   wire n_165;
   wire n_166;
   wire n_167;
   wire n_168;
   wire n_169;
   wire n_170;
   wire n_171;
   wire n_172;
   wire n_173;
   wire n_174;
   wire n_175;
   wire n_176;
   wire n_177;
   wire n_178;
   wire n_179;
   wire n_180;
   wire n_181;
   wire n_182;
   wire n_183;
   wire n_184;
   wire n_185;
   wire n_186;
   wire n_187;
   wire n_188;
   wire n_189;
   wire n_190;
   wire n_191;
   wire n_192;
   wire n_193;
   wire n_194;
   wire n_195;
   wire n_196;
   wire n_197;
   wire n_198;
   wire n_199;
   wire n_200;
   wire n_201;
   wire n_202;
   wire n_203;
   wire n_204;
   wire n_205;
   wire n_206;
   wire n_207;
   wire n_208;
   wire n_209;
   wire n_210;
   wire n_211;
   wire n_212;
   wire n_213;
   wire n_214;
   wire n_215;
   wire n_216;
   wire n_217;
   wire n_218;
   wire n_219;
   wire n_220;
   wire n_221;
   wire n_222;
   wire n_223;
   wire n_224;
   wire n_225;
   wire n_226;
   wire n_227;
   wire n_228;
   wire n_229;
   wire n_230;
   wire n_231;
   wire n_232;
   wire n_233;
   wire n_234;
   wire n_235;
   wire n_236;
   wire n_237;
   wire n_238;
   wire n_239;
   wire n_240;
   wire n_241;
   wire n_242;
   wire n_243;
   wire n_244;
   wire n_245;
   wire n_246;
   wire n_247;
   wire n_248;
   wire n_249;
   wire n_250;
   wire n_251;
   wire n_252;
   wire n_253;
   wire n_254;
   wire n_255;
   wire n_256;
   wire n_257;
   wire n_258;
   wire n_259;
   wire n_260;
   wire n_261;
   wire n_262;
   wire n_263;
   wire n_264;
   wire n_265;
   wire n_266;
   wire n_267;
   wire n_268;
   wire n_269;
   wire n_270;
   wire n_271;
   wire n_272;
   wire n_273;
   wire n_274;
   wire n_275;
   wire n_276;
   wire n_277;
   wire n_278;
   wire n_279;
   wire n_280;
   wire n_281;
   wire n_282;
   wire n_283;
   wire n_284;
   wire n_285;
   wire n_286;
   wire n_287;
   wire n_288;
   wire n_289;
   wire n_290;
   wire n_291;
   wire n_292;
   wire n_293;
   wire n_294;
   wire n_295;
   wire n_296;
   wire n_297;
   wire n_298;
   wire n_299;
   wire n_300;
   wire n_301;
   wire n_302;
   wire n_303;
   wire n_304;
   wire n_305;
   wire n_306;
   wire n_307;
   wire n_308;
   wire n_309;
   wire n_310;
   wire n_311;
   wire n_312;
   wire n_313;
   wire n_314;
   wire n_315;
   wire n_316;
   wire n_317;
   wire n_318;
   wire n_319;
   wire n_320;
   wire n_321;
   wire n_322;
   wire n_323;
   wire n_324;
   wire n_325;
   wire n_326;
   wire n_327;
   wire n_328;
   wire n_329;
   wire n_330;
   wire n_331;
   wire n_332;
   wire n_333;
   wire n_334;
   wire n_335;
   wire n_336;
   wire n_337;
   wire n_338;
   wire n_339;
   wire n_340;
   wire n_341;
   wire n_342;
   wire n_343;
   wire n_344;
   wire n_345;
   wire n_346;
   wire n_347;
   wire n_348;
   wire n_349;
   wire n_350;
   wire n_351;
   wire n_352;
   wire n_353;
   wire n_354;
   wire n_355;
   wire n_356;
   wire n_357;
   wire n_358;
   wire n_359;
   wire n_360;
   wire n_361;
   wire n_362;
   wire n_363;
   wire n_364;
   wire n_365;
   wire n_366;
   wire n_367;
   wire n_368;
   wire n_369;
   wire n_370;
   wire n_371;
   wire n_372;
   wire n_373;
   wire n_374;
   wire n_375;
   wire n_376;
   wire n_377;
   wire n_378;
   wire n_379;
   wire n_380;
   wire n_381;
   wire n_382;
   wire n_383;
   wire n_384;
   wire n_385;
   wire n_386;
   wire n_387;
   wire n_388;
   wire n_389;
   wire n_390;
   wire n_391;
   wire n_392;
   wire n_393;
   wire n_394;
   wire n_395;
   wire n_396;
   wire n_397;
   wire n_398;
   wire n_399;
   wire n_400;
   wire n_401;
   wire n_402;
   wire n_403;
   wire n_404;
   wire n_405;
   wire n_406;
   wire n_407;
   wire n_408;
   wire n_409;
   wire n_410;
   wire n_411;
   wire n_412;
   wire n_413;
   wire n_414;
   wire n_415;
   wire n_416;
   wire n_417;
   wire n_418;
   wire n_419;
   wire n_420;
   wire n_421;
   wire n_422;
   wire n_423;
   wire n_424;
   wire n_425;
   wire n_426;
   wire n_427;
   wire n_428;
   wire n_429;
   wire n_430;
   wire n_431;
   wire n_432;
   wire n_433;
   wire n_434;
   wire n_435;
   wire n_436;
   wire n_437;
   wire n_438;
   wire n_439;
   wire n_440;
   wire n_441;
   wire n_442;
   wire n_443;
   wire n_444;
   wire n_445;
   wire n_446;
   wire n_447;
   wire n_448;
   wire n_449;
   wire n_450;
   wire n_451;
   wire n_452;
   wire n_453;
   wire n_454;
   wire n_455;
   wire n_456;
   wire n_457;
   wire n_458;
   wire n_459;
   wire n_460;
   wire n_461;
   wire n_462;
   wire n_463;
   wire n_464;
   wire n_465;
   wire n_466;
   wire n_467;
   wire n_468;
   wire n_469;
   wire n_470;
   wire n_471;
   wire n_472;
   wire n_473;
   wire n_474;
   wire n_475;
   wire n_476;
   wire n_477;
   wire n_478;
   wire n_479;
   wire n_480;
   wire n_481;
   wire n_482;
   wire n_483;
   wire n_484;
   wire n_485;
   wire n_486;
   wire n_487;
   wire n_488;
   wire n_489;
   wire n_490;
   wire n_491;
   wire n_492;
   wire n_493;
   wire n_494;
   wire n_495;
   wire n_496;
   wire n_497;
   wire n_498;
   wire n_499;
   wire n_500;
   wire n_501;
   wire n_502;
   wire n_503;
   wire n_504;
   wire n_505;
   wire n_506;
   wire n_507;
   wire n_508;
   wire n_509;
   wire n_510;
   wire n_511;
   wire n_512;
   wire n_513;
   wire n_514;
   wire n_515;
   wire n_516;
   wire n_517;
   wire n_518;
   wire n_519;
   wire n_520;
   wire n_521;
   wire n_522;
   wire n_523;
   wire n_524;
   wire n_525;
   wire n_526;
   wire n_527;
   wire n_528;
   wire n_529;
   wire n_530;
   wire n_531;
   wire n_532;
   wire n_533;
   wire n_534;
   wire n_535;
   wire n_536;
   wire n_537;
   wire n_538;
   wire n_539;
   wire n_540;
   wire n_541;
   wire n_542;
   wire n_543;
   wire n_544;
   wire n_545;
   wire n_546;
   wire n_547;
   wire n_548;
   wire n_549;
   wire n_550;
   wire n_551;
   wire n_552;
   wire n_553;
   wire n_554;
   wire n_555;
   wire n_556;
   wire n_557;
   wire n_558;
   wire n_559;
   wire n_560;
   wire n_561;
   wire n_562;
   wire n_563;
   wire n_564;
   wire n_565;
   wire n_566;
   wire n_567;
   wire n_568;
   wire n_569;
   wire n_570;
   wire n_571;
   wire n_572;
   wire n_573;
   wire n_574;
   wire n_575;
   wire n_576;
   wire n_577;
   wire n_578;
   wire n_579;
   wire n_580;
   wire n_581;
   wire n_582;
   wire n_583;
   wire n_584;
   wire n_585;
   wire n_586;
   wire n_587;
   wire n_588;
   wire n_589;
   wire n_590;
   wire n_591;
   wire n_592;
   wire n_593;
   wire n_594;
   wire n_595;
   wire n_596;
   wire n_597;
   wire n_598;
   wire n_599;
   wire n_600;
   wire n_601;
   wire n_602;
   wire n_603;
   wire n_604;
   wire n_605;
   wire n_606;
   wire n_607;
   wire n_608;
   wire n_609;
   wire n_610;
   wire n_611;
   wire n_612;
   wire n_613;
   wire n_614;
   wire n_615;
   wire n_616;
   wire n_617;
   wire n_618;
   wire n_619;
   wire n_620;
   wire n_621;
   wire n_622;
   wire n_623;
   wire n_624;
   wire n_625;
   wire n_626;
   wire n_627;
   wire n_628;
   wire n_629;
   wire n_630;
   wire n_631;
   wire n_632;
   wire n_633;
   wire n_634;
   wire n_635;
   wire n_636;
   wire n_637;
   wire n_638;
   wire n_639;
   wire n_640;
   wire n_641;
   wire n_642;
   wire n_643;
   wire n_644;
   wire n_645;
   wire n_646;
   wire n_647;
   wire n_648;
   wire n_649;
   wire n_650;
   wire n_651;
   wire n_652;
   wire n_653;
   wire n_654;
   wire n_655;
   wire n_656;
   wire n_657;
   wire n_658;
   wire n_659;
   wire n_660;
   wire n_661;
   wire n_662;
   wire n_663;
   wire n_664;
   wire n_665;
   wire n_666;
   wire n_667;
   wire n_668;
   wire n_669;
   wire n_670;
   wire n_671;
   wire n_672;
   wire n_673;
   wire n_674;
   wire n_675;
   wire n_676;
   wire n_677;
   wire n_678;
   wire n_679;
   wire n_680;
   wire n_681;
   wire n_682;
   wire n_683;
   wire n_684;
   wire n_685;
   wire n_686;
   wire n_687;
   wire n_688;
   wire n_689;
   wire n_690;
   wire n_691;
   wire n_692;
   wire n_693;
   wire n_694;
   wire n_695;
   wire n_696;
   wire n_697;
   wire n_698;
   wire n_699;
   wire n_700;
   wire n_701;
   wire n_702;
   wire n_703;
   wire n_704;
   wire n_705;
   wire n_706;
   wire n_707;
   wire n_708;
   wire n_709;
   wire n_710;
   wire n_711;
   wire n_712;
   wire n_713;
   wire n_714;
   wire n_715;
   wire n_716;
   wire n_717;
   wire n_718;
   wire n_719;
   wire n_720;
   wire n_721;
   wire n_722;
   wire n_723;
   wire n_724;
   wire n_725;
   wire n_726;
   wire n_727;
   wire n_728;
   wire n_729;
   wire n_730;
   wire n_731;
   wire n_732;
   wire n_733;
   wire n_734;
   wire n_735;
   wire n_736;
   wire n_737;
   wire n_738;
   wire n_739;
   wire n_740;
   wire n_741;
   wire n_742;
   wire n_743;
   wire n_744;
   wire n_745;
   wire n_746;
   wire n_747;
   wire n_748;
   wire n_749;
   wire n_750;
   wire n_751;
   wire n_752;
   wire n_753;
   wire n_754;
   wire n_755;
   wire n_757;
   wire n_758;
   wire n_759;
   wire n_760;
   wire n_761;
   wire n_762;
   wire n_763;
   wire n_764;
   wire n_765;
   wire n_766;
   wire n_767;
   wire n_768;
   wire n_769;
   wire n_770;
   wire n_771;
   wire n_772;
   wire n_773;
   wire n_774;
   wire n_775;
   wire n_776;
   wire n_777;
   wire n_778;
   wire n_779;
   wire n_780;
   wire n_781;
   wire n_782;
   wire n_783;
   wire n_784;
   wire n_785;
   wire n_786;
   wire n_787;
   wire n_788;
   wire n_789;
   wire n_790;
   wire n_791;
   wire n_792;
   wire n_793;
   wire n_794;
   wire n_795;
   wire n_796;
   wire n_797;
   wire n_798;
   wire n_799;
   wire n_800;
   wire n_801;
   wire n_802;
   wire n_803;
   wire n_804;
   wire n_805;
   wire n_806;
   wire n_807;
   wire n_808;
   wire n_809;
   wire n_810;
   wire n_811;
   wire n_812;
   wire n_813;
   wire n_814;
   wire n_815;
   wire n_816;
   wire n_817;
   wire n_818;
   wire n_819;
   wire n_820;
   wire n_821;
   wire n_822;
   wire n_823;
   wire n_824;
   wire n_825;
   wire n_826;
   wire n_827;
   wire n_828;
   wire n_829;
   wire n_830;
   wire n_831;
   wire n_832;
   wire n_833;
   wire n_834;
   wire n_835;
   wire n_836;
   wire n_837;
   wire n_838;
   wire n_839;
   wire n_840;
   wire n_841;
   wire n_842;
   wire n_843;
   wire n_844;
   wire n_845;
   wire n_846;
   wire n_847;
   wire n_848;
   wire n_849;
   wire n_850;
   wire n_851;
   wire n_852;
   wire n_853;
   wire n_854;
   wire n_855;
   wire n_856;
   wire n_857;
   wire n_858;
   wire n_859;
   wire n_860;
   wire n_861;
   wire n_862;
   wire n_863;
   wire n_864;
   wire n_865;
   wire n_866;
   wire n_867;
   wire n_868;
   wire n_869;
   wire n_870;
   wire n_871;
   wire n_872;
   wire n_873;
   wire n_874;
   wire n_875;
   wire n_876;
   wire n_877;
   wire n_878;
   wire n_879;
   wire n_880;
   wire n_881;
   wire n_882;
   wire n_883;
   wire n_884;
   wire n_885;
   wire n_886;
   wire n_887;
   wire n_888;
   wire n_889;
   wire n_890;
   wire n_891;
   wire n_892;
   wire n_893;
   wire n_894;
   wire n_895;
   wire n_896;
   wire n_897;
   wire n_898;
   wire n_899;
   wire n_900;
   wire n_901;
   wire n_903;
   wire n_904;
   wire n_905;
   wire n_906;
   wire n_907;
   wire n_908;
   wire n_909;
   wire n_910;
   wire n_911;
   wire n_912;
   wire n_913;
   wire n_914;
   wire n_915;
   wire n_916;
   wire n_917;
   wire n_918;
   wire n_919;
   wire n_920;
   wire n_921;
   wire n_922;
   wire n_923;
   wire n_924;
   wire n_925;
   wire n_926;
   wire n_927;
   wire n_928;
   wire n_929;
   wire n_930;
   wire n_931;
   wire n_932;
   wire n_933;
   wire n_934;
   wire n_935;
   wire n_936;
   wire n_937;
   wire n_938;
   wire n_939;
   wire n_940;
   wire n_941;
   wire n_942;
   wire n_943;
   wire n_944;
   wire n_945;
   wire n_946;
   wire n_947;
   wire n_948;
   wire n_949;
   wire n_950;
   wire n_951;
   wire n_952;
   wire n_953;
   wire n_954;
   wire n_955;
   wire n_956;
   wire n_957;
   wire n_958;
   wire n_959;
   wire n_960;
   wire n_961;
   wire n_962;
   wire n_963;
   wire n_964;
   wire n_965;
   wire n_966;
   wire n_967;
   wire n_968;
   wire n_969;
   wire n_970;
   wire n_971;
   wire n_972;
   wire n_973;
   wire n_974;
   wire n_975;
   wire n_976;
   wire n_977;
   wire n_978;
   wire n_979;
   wire n_980;
   wire n_981;
   wire n_982;
   wire n_983;
   wire n_984;
   wire n_985;
   wire n_986;
   wire n_987;
   wire n_988;
   wire n_989;
   wire n_990;
   wire n_991;
   wire n_992;
   wire n_993;
   wire n_994;
   wire n_995;
   wire n_996;
   wire n_997;
   wire n_998;
   wire n_999;
   wire n_1000;
   wire n_1001;
   wire n_1002;
   wire n_1003;
   wire n_1004;
   wire n_1005;
   wire n_1006;
   wire n_1007;
   wire n_1008;
   wire n_1009;
   wire n_1011;
   wire n_1012;
   wire n_1013;
   wire n_1014;
   wire n_1015;
   wire n_1016;
   wire n_1017;
   wire n_1018;
   wire n_1019;
   wire n_1020;
   wire n_1021;
   wire n_1022;
   wire n_1023;
   wire n_1024;
   wire n_1025;
   wire n_1026;
   wire n_1027;
   wire n_1028;
   wire n_1029;
   wire n_1030;
   wire n_1031;
   wire n_1032;
   wire n_1033;
   wire n_1034;
   wire n_1035;
   wire n_1036;
   wire n_1037;
   wire n_1038;
   wire n_1039;
   wire n_1040;
   wire n_1041;
   wire n_1042;
   wire n_1043;
   wire n_1044;
   wire n_1045;
   wire n_1046;
   wire n_1047;
   wire n_1048;
   wire n_1049;
   wire n_1050;
   wire n_1051;
   wire n_1052;
   wire n_1053;
   wire n_1054;
   wire n_1055;
   wire n_1056;
   wire n_1057;
   wire n_1058;
   wire n_1059;
   wire n_1060;
   wire n_1061;
   wire n_1062;
   wire n_1063;
   wire n_1064;
   wire n_1065;
   wire n_1066;
   wire n_1067;
   wire n_1068;
   wire n_1069;
   wire n_1070;
   wire n_1071;
   wire n_1072;
   wire n_1073;
   wire n_1074;
   wire n_1075;
   wire n_1076;
   wire n_1077;
   wire n_1078;
   wire n_1079;
   wire n_1080;
   wire n_1081;
   wire n_1082;
   wire n_1083;
   wire n_1084;
   wire n_1085;
   wire n_1086;
   wire n_1087;
   wire n_1088;
   wire n_1089;
   wire n_1090;
   wire n_1091;
   wire n_1092;
   wire n_1093;
   wire n_1094;
   wire n_1095;
   wire n_1096;
   wire n_1097;
   wire n_1098;
   wire n_1099;
   wire n_1100;
   wire n_1101;
   wire n_1102;
   wire n_1103;
   wire n_1104;
   wire n_1105;
   wire n_1107;
   wire n_1108;
   wire n_1109;
   wire n_1110;
   wire n_1111;
   wire n_1112;
   wire n_1113;
   wire n_1114;
   wire n_1115;
   wire n_1116;
   wire n_1117;
   wire n_1118;
   wire n_1119;
   wire n_1120;
   wire n_1121;
   wire n_1122;
   wire n_1123;
   wire n_1124;
   wire n_1125;
   wire n_1126;
   wire n_1127;
   wire n_1128;
   wire n_1129;
   wire n_1130;
   wire n_1131;
   wire n_1132;
   wire n_1133;
   wire n_1134;
   wire n_1135;
   wire n_1136;
   wire n_1137;
   wire n_1138;
   wire n_1139;
   wire n_1140;
   wire n_1141;
   wire n_1142;
   wire n_1143;
   wire n_1144;
   wire n_1145;
   wire n_1146;
   wire n_1147;
   wire n_1148;
   wire n_1149;
   wire n_1150;
   wire n_1151;
   wire n_1152;
   wire n_1153;
   wire n_1154;
   wire n_1155;
   wire n_1156;
   wire n_1157;
   wire n_1158;
   wire n_1159;
   wire n_1160;
   wire n_1161;
   wire n_1162;
   wire n_1163;
   wire n_1164;
   wire n_1165;
   wire n_1166;
   wire n_1167;
   wire n_1168;
   wire n_1170;
   wire n_1171;
   wire n_1172;
   wire n_1173;
   wire n_1174;
   wire n_1175;
   wire n_1176;
   wire n_1177;
   wire n_1178;
   wire n_1179;
   wire n_1180;
   wire n_1181;
   wire n_1182;
   wire n_1183;
   wire n_1184;
   wire n_1185;
   wire n_1186;
   wire n_1187;
   wire n_1188;
   wire n_1189;
   wire n_1190;
   wire n_1191;
   wire n_1192;
   wire n_1193;
   wire n_1194;
   wire n_1195;
   wire n_1196;
   wire n_1197;
   wire n_1198;
   wire n_1199;
   wire n_1200;
   wire n_1201;
   wire n_1202;
   wire n_1203;
   wire n_1204;
   wire n_1205;
   wire n_1206;
   wire n_1207;
   wire n_1208;
   wire n_1209;
   wire n_1210;
   wire n_1211;
   wire n_1212;
   wire n_1213;
   wire n_1214;
   wire n_1215;
   wire n_1216;
   wire n_1217;
   wire n_1218;
   wire n_1219;
   wire n_1220;
   wire n_1221;
   wire n_1222;
   wire n_1223;
   wire n_1224;
   wire n_1225;
   wire n_1226;
   wire n_1227;
   wire n_1228;
   wire n_1229;
   wire n_1230;
   wire n_1231;
   wire n_1232;
   wire n_1233;
   wire n_1234;
   wire n_1235;
   wire n_1236;
   wire n_1237;
   wire n_1238;
   wire n_1239;
   wire n_1240;
   wire n_1242;
   wire n_1243;
   wire n_1244;
   wire n_1245;
   wire n_1246;
   wire n_1247;
   wire n_1248;
   wire n_1249;
   wire n_1250;
   wire n_1251;
   wire n_1252;
   wire n_1253;
   wire n_1254;
   wire n_1255;
   wire n_1256;
   wire n_1257;
   wire n_1258;
   wire n_1259;
   wire n_1260;
   wire n_1261;
   wire n_1262;
   wire n_1263;
   wire n_1264;
   wire n_1265;
   wire n_1266;
   wire n_1267;
   wire n_1268;
   wire n_1269;
   wire n_1270;
   wire n_1271;
   wire n_1272;
   wire n_1273;
   wire n_1274;
   wire n_1275;
   wire n_1276;
   wire n_1277;
   wire n_1278;
   wire n_1279;
   wire n_1280;
   wire n_1282;
   wire n_1283;
   wire n_1284;
   wire n_1285;
   wire n_1286;
   wire n_1287;
   wire n_1288;
   wire n_1289;
   wire n_1290;
   wire n_1291;
   wire n_1292;
   wire n_1293;
   wire n_1294;
   wire n_1295;
   wire n_1296;
   wire n_1297;
   wire n_1298;
   wire n_1299;
   wire n_1300;
   wire n_1301;
   wire n_1302;
   wire n_1303;
   wire n_1304;
   wire n_1305;
   wire n_1306;
   wire n_1307;
   wire n_1308;
   wire n_1309;
   wire n_1310;
   wire n_1311;
   wire n_1312;
   wire n_1313;
   wire n_1314;
   wire n_1315;
   wire n_1316;
   wire n_1317;
   wire n_1318;
   wire n_1320;
   wire n_1321;
   wire n_1322;
   wire n_1323;
   wire n_1324;
   wire n_1325;
   wire n_1326;
   wire n_1327;
   wire n_1328;
   wire n_1329;
   wire n_1330;
   wire n_1331;
   wire n_1332;
   wire n_1333;
   wire n_1334;
   wire n_1335;
   wire n_1336;
   wire n_1337;
   wire n_1339;
   wire n_1340;
   wire n_1341;
   wire n_1342;
   wire n_1343;
   wire n_1344;
   wire n_1345;
   wire n_1346;
   wire n_1347;
   wire n_1348;
   wire n_1349;
   wire n_1350;
   wire n_1351;
   wire n_1352;
   wire n_1353;
   wire n_1354;
   wire n_1356;
   wire n_1357;
   wire n_1358;
   wire n_1359;
   wire n_1361;
   wire n_1362;
   wire n_1364;
   wire n_1365;
   wire n_1367;
   wire n_1368;
   wire n_1370;
   wire n_1371;
   wire n_1373;
   wire n_1374;
   wire n_1376;
   wire n_1377;
   wire n_1379;
   wire n_1380;
   wire n_1382;
   wire n_1383;
   wire n_1385;
   wire n_1386;
   wire n_1388;
   wire n_1389;
   wire n_1391;
   wire n_1392;
   wire n_1394;
   wire n_1395;
   wire n_1397;
   wire n_1398;
   wire n_1400;
   wire n_1401;
   wire n_1403;
   wire n_1404;
   wire n_1406;
   wire n_1407;
   wire n_1409;
   wire n_1410;
   wire n_1412;
   wire n_1413;
   wire n_1415;
   wire n_1416;
   wire n_1418;
   wire n_1419;
   wire n_1421;
   wire n_1422;
   wire n_1424;
   wire n_1425;
   wire n_1427;
   wire n_1428;
   wire n_1430;
   wire n_1431;
   wire n_1433;
   wire n_1434;
   wire n_1436;
   wire n_1437;
   wire n_1439;
   wire n_1440;
   wire n_1442;
   wire n_1443;
   wire n_1445;
   wire n_1446;
   wire n_1448;
   wire n_1449;
   wire n_1451;
   wire n_1452;
   wire n_1454;
   wire n_1455;
   wire n_1457;
   wire n_1458;
   wire n_1460;
   wire n_1461;
   wire n_1463;
   wire n_1464;

   EN3X1 g28144 (.Q(Z[47]), 
	.C(n_1463), 
	.B(n_999), 
	.A(n_792));
   INX4 g28145 (.Q(Z[46]), 
	.A(n_1464));
   FAX4 g28146 (.S(n_1464), 
	.CO(n_1463), 
	.CI(n_1460), 
	.B(n_1029), 
	.A(n_1000));
   INX4 g28147 (.Q(Z[45]), 
	.A(n_1461));
   FAX4 g28148 (.S(n_1461), 
	.CO(n_1460), 
	.CI(n_1457), 
	.B(n_1030), 
	.A(n_1142));
   INX4 g28149 (.Q(Z[44]), 
	.A(n_1458));
   FAX4 g28150 (.S(n_1458), 
	.CO(n_1457), 
	.CI(n_1454), 
	.B(n_1182), 
	.A(n_1143));
   INX4 g28151 (.Q(Z[43]), 
	.A(n_1455));
   FAX4 g28152 (.S(n_1455), 
	.CO(n_1454), 
	.CI(n_1451), 
	.B(n_1248), 
	.A(n_1183));
   INX4 g28153 (.Q(Z[42]), 
	.A(n_1452));
   FAX4 g28154 (.S(n_1452), 
	.CO(n_1451), 
	.CI(n_1448), 
	.B(n_1249), 
	.A(n_1204));
   INX4 g28155 (.Q(Z[41]), 
	.A(n_1449));
   FAX4 g28156 (.S(n_1449), 
	.CO(n_1448), 
	.CI(n_1445), 
	.B(n_1205), 
	.A(n_1242));
   INX4 g28157 (.Q(Z[40]), 
	.A(n_1446));
   FAX4 g28158 (.S(n_1446), 
	.CO(n_1445), 
	.CI(n_1442), 
	.B(n_1285), 
	.A(n_1243));
   INX4 g28159 (.Q(Z[39]), 
	.A(n_1443));
   FAX4 g28160 (.S(n_1443), 
	.CO(n_1442), 
	.CI(n_1439), 
	.B(n_1286), 
	.A(n_1275));
   INX4 g28161 (.Q(Z[38]), 
	.A(n_1440));
   FAX4 g28162 (.S(n_1440), 
	.CO(n_1439), 
	.CI(n_1436), 
	.B(n_1276), 
	.A(n_1292));
   INX4 g28163 (.Q(Z[37]), 
	.A(n_1437));
   FAX4 g28164 (.S(n_1437), 
	.CO(n_1436), 
	.CI(n_1433), 
	.B(n_1313), 
	.A(n_1293));
   INX4 g28165 (.Q(Z[36]), 
	.A(n_1434));
   FAX4 g28166 (.S(n_1434), 
	.CO(n_1433), 
	.CI(n_1430), 
	.B(n_1314), 
	.A(n_1328));
   INX4 g28167 (.Q(Z[35]), 
	.A(n_1431));
   FAX4 g28168 (.S(n_1431), 
	.CO(n_1430), 
	.CI(n_1427), 
	.B(n_1329), 
	.A(n_1322));
   INX4 g28169 (.Q(Z[34]), 
	.A(n_1428));
   FAX4 g28170 (.S(n_1428), 
	.CO(n_1427), 
	.CI(n_1424), 
	.B(n_11), 
	.A(n_1325));
   INX4 g28171 (.Q(Z[33]), 
	.A(n_1425));
   FAX4 g28172 (.S(n_1425), 
	.CO(n_1424), 
	.CI(n_1421), 
	.B(n_1326), 
	.A(n_1327));
   INX4 g28173 (.Q(Z[32]), 
	.A(n_1422));
   FAX4 g28174 (.S(n_1422), 
	.CO(n_1421), 
	.CI(n_1418), 
	.B(n_12), 
	.A(n_1339));
   INX4 g28175 (.Q(Z[31]), 
	.A(n_1419));
   FAX4 g28176 (.S(n_1419), 
	.CO(n_1418), 
	.CI(n_1415), 
	.B(n_1340), 
	.A(n_1356));
   INX4 g28177 (.Q(Z[30]), 
	.A(n_1416));
   FAX4 g28178 (.S(n_1416), 
	.CO(n_1415), 
	.CI(n_1412), 
	.B(n_1351), 
	.A(n_1357));
   INX4 g28179 (.Q(Z[29]), 
	.A(n_1413));
   FAX4 g28180 (.S(n_1413), 
	.CO(n_1412), 
	.CI(n_1409), 
	.B(n_1352), 
	.A(n_1349));
   INX4 g28181 (.Q(Z[28]), 
	.A(n_1410));
   FAX4 g28182 (.S(n_1410), 
	.CO(n_1409), 
	.CI(n_1406), 
	.B(n_1350), 
	.A(n_1347));
   INX4 g28183 (.Q(Z[27]), 
	.A(n_1407));
   FAX4 g28184 (.S(n_1407), 
	.CO(n_1406), 
	.CI(n_1403), 
	.B(n_1345), 
	.A(n_1348));
   INX4 g28185 (.Q(Z[26]), 
	.A(n_1404));
   FAX4 g28186 (.S(n_1404), 
	.CO(n_1403), 
	.CI(n_1400), 
	.B(n_1346), 
	.A(n_1343));
   INX4 g28187 (.Q(Z[25]), 
	.A(n_1401));
   FAX4 g28188 (.S(n_1401), 
	.CO(n_1400), 
	.CI(n_1397), 
	.B(n_1344), 
	.A(n_1341));
   INX4 g28189 (.Q(Z[24]), 
	.A(n_1398));
   FAX4 g28190 (.S(n_1398), 
	.CO(n_1397), 
	.CI(n_1394), 
	.B(n_1342), 
	.A(n_1332));
   INX4 g28191 (.Q(Z[23]), 
	.A(n_1395));
   FAX4 g28192 (.S(n_1395), 
	.CO(n_1394), 
	.CI(n_1391), 
	.B(n_1333), 
	.A(n_1330));
   INX4 g28193 (.Q(Z[22]), 
	.A(n_1392));
   FAX4 g28194 (.S(n_1392), 
	.CO(n_1391), 
	.CI(n_1388), 
	.B(n_1331), 
	.A(n_1334));
   INX4 g28195 (.Q(Z[21]), 
	.A(n_1389));
   FAX4 g28196 (.S(n_1389), 
	.CO(n_1388), 
	.CI(n_1385), 
	.B(n_1335), 
	.A(n_1309));
   INX4 g28197 (.Q(Z[20]), 
	.A(n_1386));
   FAX4 g28198 (.S(n_1386), 
	.CO(n_1385), 
	.CI(n_1382), 
	.B(n_1305), 
	.A(n_1310));
   INX4 g28199 (.Q(Z[19]), 
	.A(n_1383));
   FAX4 g28200 (.S(n_1383), 
	.CO(n_1382), 
	.CI(n_1379), 
	.B(n_1306), 
	.A(n_1301));
   INX4 g28201 (.Q(Z[18]), 
	.A(n_1380));
   FAX4 g28202 (.S(n_1380), 
	.CO(n_1379), 
	.CI(n_1376), 
	.B(n_1299), 
	.A(n_1302));
   INX4 g28203 (.Q(Z[17]), 
	.A(n_1377));
   FAX4 g28204 (.S(n_1377), 
	.CO(n_1376), 
	.CI(n_1373), 
	.B(n_1300), 
	.A(n_1277));
   INX4 g28205 (.Q(Z[16]), 
	.A(n_1374));
   FAX4 g28206 (.S(n_1374), 
	.CO(n_1373), 
	.CI(n_1370), 
	.B(n_1278), 
	.A(n_1265));
   INX4 g28207 (.Q(Z[15]), 
	.A(n_1371));
   FAX4 g28208 (.S(n_1371), 
	.CO(n_1370), 
	.CI(n_1367), 
	.B(n_1266), 
	.A(n_1283));
   INX4 g28209 (.Q(Z[14]), 
	.A(n_1368));
   FAX4 g28210 (.S(n_1368), 
	.CO(n_1367), 
	.CI(n_1364), 
	.B(n_1284), 
	.A(n_1210));
   INX4 g28211 (.Q(Z[13]), 
	.A(n_1365));
   FAX4 g28212 (.S(n_1365), 
	.CO(n_1364), 
	.CI(n_1361), 
	.B(n_1192), 
	.A(n_1211));
   INX4 g28213 (.Q(Z[12]), 
	.A(n_1362));
   FAX4 g28214 (.S(n_1362), 
	.CO(n_1361), 
	.CI(n_1358), 
	.B(n_1193), 
	.A(n_1190));
   INX4 g28215 (.Q(Z[11]), 
	.A(n_1359));
   FAX4 g28216 (.S(n_1359), 
	.CO(n_1358), 
	.CI(n_1353), 
	.B(n_1191), 
	.A(n_1161));
   FAX4 g28217 (.S(n_1357), 
	.CO(n_1356), 
	.CI(n_1303), 
	.B(n_1308), 
	.A(n_1253));
   INX4 g28218 (.Q(Z[10]), 
	.A(n_1354));
   FAX4 g28219 (.S(n_1354), 
	.CO(n_1353), 
	.CI(n_1336), 
	.B(n_1162), 
	.A(n_1113));
   FAX4 g28220 (.S(n_1352), 
	.CO(n_1351), 
	.CI(n_1304), 
	.B(n_1295), 
	.A(n_1206));
   FAX4 g28221 (.S(n_1350), 
	.CO(n_1349), 
	.CI(n_1320), 
	.B(n_1296), 
	.A(n_1207));
   FAX4 g28222 (.S(n_1348), 
	.CO(n_1347), 
	.CI(n_1321), 
	.B(n_1315), 
	.A(n_1209));
   FAX4 g28223 (.S(n_1346), 
	.CO(n_1345), 
	.CI(n_1316), 
	.B(n_1311), 
	.A(n_1257));
   FAX4 g28224 (.S(n_1344), 
	.CO(n_1343), 
	.CI(n_1312), 
	.B(n_1297), 
	.A(n_1229));
   FAX4 g28225 (.S(n_1342), 
	.CO(n_1341), 
	.CI(n_1290), 
	.B(n_1298), 
	.A(n_1230));
   FAX4 g28226 (.S(n_1340), 
	.CO(n_1339), 
	.CI(n_1307), 
	.B(n_1287), 
	.A(n_1228));
   INX4 g28227 (.Q(Z[9]), 
	.A(n_1337));
   FAX4 g28228 (.S(n_1337), 
	.CO(n_1336), 
	.CI(n_1317), 
	.B(n_1114), 
	.A(n_1023));
   FAX4 g28229 (.S(n_1335), 
	.CO(n_1334), 
	.CI(n_1270), 
	.B(n_1267), 
	.A(n_1216));
   FAX4 g28230 (.S(n_1333), 
	.CO(n_1332), 
	.CI(n_1291), 
	.B(n_1271), 
	.A(n_1222));
   FAX4 g28231 (.S(n_1331), 
	.CO(n_1330), 
	.CI(n_1269), 
	.B(n_1272), 
	.A(n_1223));
   FAX4 g28233 (.S(n_1329), 
	.CO(n_1328), 
	.CI(n_1258), 
	.B(n_1262), 
	.A(n_1118));
   EN3X2 g28235 (.Q(n_1327), 
	.C(n_1289), 
	.B(n_1274), 
	.A(n_1203));
   INX8789 g28237 (.Q(n_1326), 
	.A(n_1324));
   INX8 g28238 (.Q(n_1325), 
	.A(n_1323));
   FAX3 g28239 (.S(n_1324), 
	.CO(n_1323), 
	.CI(n_1263), 
	.B(n_1254), 
	.A(n_1273));
   EN3X2 g28240 (.Q(n_1322), 
	.C(n_1264), 
	.B(n_1260), 
	.A(n_1255));
   FAX4 g28242 (.S(n_1321), 
	.CO(n_1320), 
	.CI(n_1195), 
	.B(n_1235), 
	.A(n_1256));
   INX4 g28243 (.Q(Z[8]), 
	.A(n_1318));
   FAX4 g28244 (.S(n_1318), 
	.CO(n_1317), 
	.CI(n_1279), 
	.B(n_1024), 
	.A(n_1045));
   FAX3 g28245 (.S(n_1316), 
	.CO(n_1315), 
	.CI(n_1231), 
	.B(n_1233), 
	.A(n_1236));
   FAX4 g28246 (.S(n_1314), 
	.CO(n_1313), 
	.CI(n_1199), 
	.B(n_1261), 
	.A(n_1117));
   FAX3 g28247 (.S(n_1312), 
	.CO(n_1311), 
	.CI(n_1234), 
	.B(n_1200), 
	.A(n_1232));
   FAX4 g28248 (.S(n_1310), 
	.CO(n_1309), 
	.CI(n_1268), 
	.B(n_1196), 
	.A(n_1184));
   FAX4 g28249 (.S(n_1308), 
	.CO(n_1307), 
	.CI(n_1218), 
	.B(n_1214), 
	.A(n_1166));
   FAX4 g28250 (.S(n_1306), 
	.CO(n_1305), 
	.CI(n_1197), 
	.B(n_1244), 
	.A(n_1185));
   FAX3 g28251 (.S(n_1304), 
	.CO(n_1303), 
	.CI(n_1219), 
	.B(n_1160), 
	.A(n_1215));
   FAX4 g28252 (.S(n_1302), 
	.CO(n_1301), 
	.CI(n_1245), 
	.B(n_1212), 
	.A(n_1130));
   FAX4 g28253 (.S(n_1300), 
	.CO(n_1299), 
	.CI(n_1213), 
	.B(n_1237), 
	.A(n_1070));
   FAX4 g28254 (.S(n_1298), 
	.CO(n_1297), 
	.CI(n_1224), 
	.B(n_1201), 
	.A(n_1188));
   FAX4 g28255 (.S(n_1296), 
	.CO(n_1295), 
	.CI(n_1208), 
	.B(n_10), 
	.A(n_1194));
   EO2X3 g28256 (.Q(n_1294), 
	.B(n_1274), 
	.A(n_1203));
   FAX4 g28257 (.S(n_1293), 
	.CO(n_1292), 
	.CI(n_1198), 
	.B(n_1187), 
	.A(n_1108));
   FAX3 g28258 (.S(n_1291), 
	.CO(n_1290), 
	.CI(n_1225), 
	.B(n_1138), 
	.A(n_1189));
   INCX4 g28259 (.Q(n_1289), 
	.A(n_1288));
   FAX4 g28260 (.S(n_1287), 
	.CO(n_1288), 
	.CI(n_1252), 
	.B(n_1151), 
	.A(n_1165));
   FAX4 g28261 (.S(n_1286), 
	.CO(n_1285), 
	.CI(n_1170), 
	.B(n_1179), 
	.A(n_1056));
   FAX4 g28262 (.S(n_1284), 
	.CO(n_1283), 
	.CI(n_1173), 
	.B(n_1121), 
	.A(n_1059));
   EN2X4 g28263 (.Q(n_1282), 
	.B(n_1259), 
	.A(n_1255));
   INX4 g28264 (.Q(Z[7]), 
	.A(n_1280));
   FAX4 g28265 (.S(n_1280), 
	.CO(n_1279), 
	.CI(n_1239), 
	.B(n_1046), 
	.A(n_993));
   FAX4 g28266 (.S(n_1278), 
	.CO(n_1277), 
	.CI(n_1238), 
	.B(n_1068), 
	.A(n_1163));
   FAX4 g28267 (.S(n_1276), 
	.CO(n_1275), 
	.CI(n_1186), 
	.B(n_1171), 
	.A(n_1057));
   FAX4 g28268 (.S(n_1274), 
	.CO(n_1273), 
	.CI(n_1226), 
	.B(n_1103), 
	.A(n_1152));
   FAX4 g28269 (.S(n_1272), 
	.CO(n_1271), 
	.CI(n_1220), 
	.B(n_1091), 
	.A(n_1139));
   FAX3 g28270 (.S(n_1270), 
	.CO(n_1269), 
	.CI(n_1221), 
	.B(n_1082), 
	.A(n_1089));
   FAX3 g28271 (.S(n_1268), 
	.CO(n_1267), 
	.CI(n_1217), 
	.B(n_1132), 
	.A(n_1083));
   FAX4 g28272 (.S(n_1266), 
	.CO(n_1265), 
	.CI(n_1164), 
	.B(n_1052), 
	.A(n_1172));
   FAX3 g28273 (.S(n_1263), 
	.CO(n_1264), 
	.CI(n_1202), 
	.B(n_1102), 
	.A(n_1055));
   FAX4 g28274 (.S(n_1262), 
	.CO(n_1261), 
	.CI(n_1176), 
	.B(n_1032), 
	.A(n_1063));
   INX8 g28275 (.Q(n_1260), 
	.A(n_1259));
   FAX4 g28276 (.S(n_1259), 
	.CO(n_1258), 
	.CI(n_1177), 
	.B(n_1053), 
	.A(n_1064));
   FAX4 g28277 (.S(n_1257), 
	.CO(n_1256), 
	.CI(n_1043), 
	.B(n_1042), 
	.A(n_1155));
   FAX4 g28278 (.S(n_1254), 
	.CO(n_1255), 
	.CI(n_1072), 
	.B(n_1157), 
	.A(n_962));
   INX8 g28279 (.Q(n_1253), 
	.A(n_1251));
   INX8 g28280 (.Q(n_1252), 
	.A(n_1250));
   FAX4 g28281 (.S(n_1251), 
	.CO(n_1250), 
	.CI(n_1093), 
	.B(n_1149), 
	.A(n_1133));
   INX8 g28282 (.Q(n_1249), 
	.A(n_1247));
   INX8 g28283 (.Q(n_1248), 
	.A(n_1246));
   FAX3 g28284 (.S(n_1247), 
	.CO(n_1246), 
	.CI(n_1011), 
	.B(n_933), 
	.A(n_1145));
   FAX3 g28285 (.S(n_1245), 
	.CO(n_1244), 
	.CI(n_1078), 
	.B(n_1125), 
	.A(n_1069));
   FAX4 g28286 (.S(n_1243), 
	.CO(n_1242), 
	.CI(n_1178), 
	.B(n_1154), 
	.A(n_1136));
   INX4 g28287 (.Q(Z[6]), 
	.A(n_1240));
   FAX4 g28288 (.S(n_1240), 
	.CO(n_1239), 
	.CI(n_1167), 
	.B(n_994), 
	.A(n_986));
   FAX3 g28289 (.S(n_1238), 
	.CO(n_1237), 
	.CI(n_1051), 
	.B(n_1001), 
	.A(n_1066));
   FAX4 g28290 (.S(n_1236), 
	.CO(n_1235), 
	.CI(n_1116), 
	.B(n_1109), 
	.A(n_1050));
   FAX3 g28291 (.S(n_1234), 
	.CO(n_1233), 
	.CI(n_1100), 
	.B(n_1020), 
	.A(n_1110));
   FAX4 g28292 (.S(n_1232), 
	.CO(n_1231), 
	.CI(n_1044), 
	.B(n_1037), 
	.A(n_1156));
   FAX4 g28293 (.S(n_1230), 
	.CO(n_1229), 
	.CI(n_1038), 
	.B(n_1094), 
	.A(n_1101));
   INX8 g28294 (.Q(n_1228), 
	.A(n_1227));
   FAX4 g28295 (.S(n_1227), 
	.CO(n_1226), 
	.CI(n_1092), 
	.B(n_1099), 
	.A(n_1148));
   FAX3 g28296 (.S(n_1225), 
	.CO(n_1224), 
	.CI(n_1095), 
	.B(n_1097), 
	.A(n_1090));
   FAX3 g28297 (.S(n_1223), 
	.CO(n_1222), 
	.CI(n_1088), 
	.B(n_1084), 
	.A(n_1147));
   FAX3 g28298 (.S(n_1221), 
	.CO(n_1220), 
	.CI(n_1085), 
	.B(n_1131), 
	.A(n_1019));
   FAX3 g28299 (.S(n_1219), 
	.CO(n_1218), 
	.CI(n_1135), 
	.B(n_1087), 
	.A(n_1127));
   FAX3 g28300 (.S(n_1217), 
	.CO(n_1216), 
	.CI(n_1075), 
	.B(n_8), 
	.A(n_1073));
   FAX4 g28301 (.S(n_1215), 
	.CO(n_1214), 
	.CI(n_1080), 
	.B(n_1005), 
	.A(n_863));
   FAX3 g28302 (.S(n_1213), 
	.CO(n_1212), 
	.CI(n_1067), 
	.B(n_1065), 
	.A(n_1126));
   FAX4 g28303 (.S(n_1211), 
	.CO(n_1210), 
	.CI(n_1122), 
	.B(n_1119), 
	.A(n_1124));
   FAX4 g28304 (.S(n_1209), 
	.CO(n_1208), 
	.CI(n_1112), 
	.B(n_1048), 
	.A(n_1115));
   FAX4 g28305 (.S(n_1207), 
	.CO(n_1206), 
	.CI(n_1128), 
	.B(n_1111), 
	.A(n_1047));
   FAX4 g28306 (.S(n_1205), 
	.CO(n_1204), 
	.CI(n_1022), 
	.B(n_1153), 
	.A(n_1003));
   FAX4 g28307 (.S(n_1203), 
	.CO(n_1202), 
	.CI(n_1158), 
	.B(n_1098), 
	.A(n_991));
   FAX3 g28308 (.S(n_1201), 
	.CO(n_1200), 
	.CI(n_1096), 
	.B(n_964), 
	.A(n_1021));
   FAX3 g28309 (.S(n_1199), 
	.CO(n_1198), 
	.CI(n_1040), 
	.B(n_1036), 
	.A(n_1031));
   FAX4 g28310 (.S(n_1197), 
	.CO(n_1196), 
	.CI(n_1076), 
	.B(n_1129), 
	.A(n_1077));
   FAX3 g28312 (.S(n_1195), 
	.CO(n_1194), 
	.CI(n_1041), 
	.B(n_1049), 
	.A(n_1062));
   FAX4 g28313 (.S(n_1193), 
	.CO(n_1192), 
	.CI(n_1120), 
	.B(n_1025), 
	.A(n_1017));
   FAX4 g28314 (.S(n_1191), 
	.CO(n_1190), 
	.CI(n_1033), 
	.B(n_1026), 
	.A(n_971));
   FAX4 g28315 (.S(n_1189), 
	.CO(n_1188), 
	.CI(n_1146), 
	.B(n_965), 
	.A(n_893));
   FAX4 g28316 (.S(n_1187), 
	.CO(n_1186), 
	.CI(n_1039), 
	.B(n_1035), 
	.A(n_996));
   FAX4 g28317 (.S(n_1185), 
	.CO(n_1184), 
	.CI(n_1074), 
	.B(n_997), 
	.A(n_936));
   INX8 g28318 (.Q(n_1183), 
	.A(n_1181));
   INX8 g28319 (.Q(n_1182), 
	.A(n_1180));
   FAX3 g28320 (.S(n_1181), 
	.CO(n_1180), 
	.CI(n_1144), 
	.B(n_845), 
	.A(n_1015));
   FAX4 g28321 (.S(n_1179), 
	.CO(n_1178), 
	.CI(n_1137), 
	.B(n_891), 
	.A(n_786));
   INX8 g28322 (.Q(n_1177), 
	.A(n_1175));
   INX8 g28323 (.Q(n_1176), 
	.A(n_1174));
   FAX3 g28324 (.S(n_1175), 
	.CO(n_1174), 
	.CI(n_1071), 
	.B(n_791), 
	.A(n_989));
   FAX3 g28325 (.S(n_1173), 
	.CO(n_1172), 
	.CI(n_1123), 
	.B(n_7), 
	.A(n_828));
   FAX4 g28327 (.S(n_1171), 
	.CO(n_1170), 
	.CI(n_1107), 
	.B(n_995), 
	.A(n_4));
   INX4 g28328 (.Q(Z[5]), 
	.A(n_1168));
   FAX4 g28329 (.S(n_1168), 
	.CO(n_1167), 
	.CI(n_1104), 
	.B(n_987), 
	.A(n_856));
   FAX4 g28330 (.S(n_1166), 
	.CO(n_1165), 
	.CI(n_1086), 
	.B(n_796), 
	.A(n_862));
   FAX3 g28331 (.S(n_1164), 
	.CO(n_1163), 
	.CI(n_1058), 
	.B(n_793), 
	.A(n_1002));
   FAX4 g28332 (.S(n_1162), 
	.CO(n_1161), 
	.CI(n_1034), 
	.B(n_1012), 
	.A(n_869));
   EN3X2 g28333 (.Q(n_1160), 
	.C(n_1081), 
	.B(n_1061), 
	.A(n_1007));
   EN2X4 g28334 (.Q(n_1159), 
	.B(n_1061), 
	.A(n_1007));
   FAX3 g28335 (.S(n_1158), 
	.CO(n_1157), 
	.CI(n_809), 
	.B(n_799), 
	.A(n_911));
   FAX3 g28336 (.S(n_1156), 
	.CO(n_1155), 
	.CI(n_982), 
	.B(n_874), 
	.A(n_788));
   FAX4 g28337 (.S(n_1154), 
	.CO(n_1153), 
	.CI(n_1004), 
	.B(n_789), 
	.A(n_890));
   INX8 g28338 (.Q(n_1152), 
	.A(n_1150));
   FAX4 g28339 (.S(n_1151), 
	.CO(n_1150), 
	.CI(n_990), 
	.B(n_800), 
	.A(n_806));
   FAX4 g28340 (.S(n_1149), 
	.CO(n_1148), 
	.CI(n_958), 
	.B(n_954), 
	.A(n_692));
   FAX4 g28341 (.S(n_1147), 
	.CO(n_1146), 
	.CI(n_948), 
	.B(n_872), 
	.A(n_758));
   FAX4 g28342 (.S(n_1145), 
	.CO(n_1144), 
	.CI(n_920), 
	.B(n_950), 
	.A(n_693));
   INX8 g28343 (.Q(n_1143), 
	.A(n_1141));
   INX8 g28344 (.Q(n_1142), 
	.A(n_1140));
   FAX3 g28345 (.S(n_1141), 
	.CO(n_1140), 
	.CI(n_1014), 
	.B(n_844), 
	.A(n_851));
   FAX4 g28346 (.S(n_1139), 
	.CO(n_1138), 
	.CI(n_1018), 
	.B(n_916), 
	.A(n_904));
   FAX3 g28347 (.S(n_1137), 
	.CO(n_1136), 
	.CI(n_879), 
	.B(n_528), 
	.A(n_941));
   INX8 g28348 (.Q(n_1135), 
	.A(n_1134));
   FAX3 g28349 (.S(n_1134), 
	.CO(n_1133), 
	.CI(n_959), 
	.B(n_947), 
	.A(n_955));
   FAX4 g28350 (.S(n_1132), 
	.CO(n_1131), 
	.CI(n_935), 
	.B(n_923), 
	.A(n_882));
   FAX4 g28351 (.S(n_1130), 
	.CO(n_1129), 
	.CI(n_998), 
	.B(n_937), 
	.A(n_855));
   FAX4 g28352 (.S(n_1128), 
	.CO(n_1127), 
	.CI(n_940), 
	.B(n_914), 
	.A(n_861));
   FAX3 g28353 (.S(n_1126), 
	.CO(n_1125), 
	.CI(n_976), 
	.B(n_880), 
	.A(n_956));
   FAX3 g28354 (.S(n_1124), 
	.CO(n_1123), 
	.CI(n_925), 
	.B(n_749), 
	.A(n_978));
   FAX4 g28355 (.S(n_1122), 
	.CO(n_1121), 
	.CI(n_1016), 
	.B(n_985), 
	.A(n_930));
   FAX3 g28356 (.S(n_1120), 
	.CO(n_1119), 
	.CI(n_970), 
	.B(n_979), 
	.A(n_926));
   FAX4 g28357 (.S(n_1118), 
	.CO(n_1117), 
	.CI(n_988), 
	.B(n_9), 
	.A(n_843));
   FAX3 g28358 (.S(n_1116), 
	.CO(n_1115), 
	.CI(n_797), 
	.B(n_967), 
	.A(n_830));
   FAX4 g28359 (.S(n_1114), 
	.CO(n_1113), 
	.CI(n_1013), 
	.B(n_818), 
	.A(n_795));
   FAX3 g28360 (.S(n_1112), 
	.CO(n_1111), 
	.CI(n_801), 
	.B(n_829), 
	.A(n_798));
   FAX4 g28361 (.S(n_1110), 
	.CO(n_1109), 
	.CI(n_906), 
	.B(n_968), 
	.A(n_676));
   FAX4 g28362 (.S(n_1108), 
	.CO(n_1107), 
	.CI(n_918), 
	.B(n_922), 
	.A(n_858));
   INX4 g28363 (.Q(Z[4]), 
	.A(n_1105));
   FAX4 g28364 (.S(n_1105), 
	.CO(n_1104), 
	.CI(n_1008), 
	.B(n_857), 
	.A(n_747));
   FAX3 g28365 (.S(n_1103), 
	.CO(n_1102), 
	.CI(n_928), 
	.B(n_963), 
	.A(n_839));
   FAX4 g28366 (.S(n_1101), 
	.CO(n_1100), 
	.CI(n_969), 
	.B(n_892), 
	.A(n_974));
   FAX4 g28367 (.S(n_1099), 
	.CO(n_1098), 
	.CI(n_912), 
	.B(n_972), 
	.A(n_805));
   FAX4 g28368 (.S(n_1097), 
	.CO(n_1096), 
	.CI(n_960), 
	.B(n_915), 
	.A(n_903));
   FAX3 g28369 (.S(n_1095), 
	.CO(n_1094), 
	.CI(n_975), 
	.B(n_952), 
	.A(n_849));
   FAX3 g28370 (.S(n_1093), 
	.CO(n_1092), 
	.CI(n_810), 
	.B(n_946), 
	.A(n_973));
   FAX4 g28371 (.S(n_1091), 
	.CO(n_1090), 
	.CI(n_961), 
	.B(n_953), 
	.A(n_870));
   FAX3 g28372 (.S(n_1089), 
	.CO(n_1088), 
	.CI(n_873), 
	.B(n_794), 
	.A(n_871));
   FAX4 g28373 (.S(n_1087), 
	.CO(n_1086), 
	.CI(n_939), 
	.B(n_913), 
	.A(n_860));
   FAX3 g28374 (.S(n_1085), 
	.CO(n_1084), 
	.CI(n_949), 
	.B(n_815), 
	.A(n_825));
   FAX4 g28375 (.S(n_1083), 
	.CO(n_1082), 
	.CI(n_826), 
	.B(n_865), 
	.A(n_816));
   INX8 g28376 (.Q(n_1080), 
	.A(n_1079));
   FAX4 g28377 (.S(n_1081), 
	.CO(n_1079), 
	.CI(n_808), 
	.B(n_943), 
	.A(n_804));
   FAX3 g28378 (.S(n_1078), 
	.CO(n_1077), 
	.CI(n_932), 
	.B(n_885), 
	.A(n_846));
   FAX4 g28379 (.S(n_1076), 
	.CO(n_1075), 
	.CI(n_924), 
	.B(n_883), 
	.A(n_931));
   FAX4 g28380 (.S(n_1074), 
	.CO(n_1073), 
	.CI(n_854), 
	.B(n_884), 
	.A(n_752));
   FAX4 g28381 (.S(n_1072), 
	.CO(n_1071), 
	.CI(n_927), 
	.B(n_838), 
	.A(n_702));
   FAX4 g28382 (.S(n_1070), 
	.CO(n_1069), 
	.CI(n_847), 
	.B(n_938), 
	.A(n_853));
   FAX4 g28383 (.S(n_1068), 
	.CO(n_1067), 
	.CI(n_977), 
	.B(n_957), 
	.A(n_881));
   FAX4 g28384 (.S(n_1066), 
	.CO(n_1065), 
	.CI(n_980), 
	.B(n_907), 
	.A(n_741));
   FAX4 g28385 (.S(n_1064), 
	.CO(n_1063), 
	.CI(n_867), 
	.B(n_888), 
	.A(n_831));
   INX8 g28386 (.Q(n_1062), 
	.A(n_1060));
   FAX3 g28387 (.S(n_1060), 
	.CO(n_1061), 
	.CI(n_803), 
	.B(n_558), 
	.A(n_833));
   FAX4 g28388 (.S(n_1059), 
	.CO(n_1058), 
	.CI(n_984), 
	.B(n_929), 
	.A(n_887));
   FAX4 g28389 (.S(n_1057), 
	.CO(n_1056), 
	.CI(n_942), 
	.B(n_921), 
	.A(n_917));
   INX8 g28390 (.Q(n_1055), 
	.A(n_1054));
   FAX3 g28391 (.S(n_1054), 
	.CO(n_1053), 
	.CI(n_802), 
	.B(n_832), 
	.A(n_889));
   FAX3 g28392 (.S(n_1052), 
	.CO(n_1051), 
	.CI(n_981), 
	.B(n_827), 
	.A(n_908));
   FAX4 g28393 (.S(n_1050), 
	.CO(n_1049), 
	.CI(n_905), 
	.B(n_896), 
	.A(n_819));
   FAX4 g28394 (.S(n_1048), 
	.CO(n_1047), 
	.CI(n_945), 
	.B(n_837), 
	.A(n_966));
   FAX4 g28395 (.S(n_1046), 
	.CO(n_1045), 
	.CI(n_910), 
	.B(n_813), 
	.A(n_755));
   FAX3 g28396 (.S(n_1044), 
	.CO(n_1043), 
	.CI(n_895), 
	.B(n_820), 
	.A(n_897));
   FAX4 g28397 (.S(n_1042), 
	.CO(n_1041), 
	.CI(n_835), 
	.B(n_894), 
	.A(n_677));
   FAX3 g28398 (.S(n_1040), 
	.CO(n_1039), 
	.CI(n_859), 
	.B(n_842), 
	.A(n_824));
   FAX4 g28399 (.S(n_1038), 
	.CO(n_1037), 
	.CI(n_5), 
	.B(n_983), 
	.A(n_875));
   FAX4 g28400 (.S(n_1036), 
	.CO(n_1035), 
	.CI(n_821), 
	.B(n_812), 
	.A(n_695));
   FAX4 g28401 (.S(n_1034), 
	.CO(n_1033), 
	.CI(n_841), 
	.B(n_817), 
	.A(n_759));
   FAX4 g28402 (.S(n_1032), 
	.CO(n_1031), 
	.CI(n_822), 
	.B(n_787), 
	.A(n_866));
   INX8 g28403 (.Q(n_1030), 
	.A(n_1028));
   INX8 g28404 (.Q(n_1029), 
	.A(n_1027));
   FAX3 g28405 (.S(n_1028), 
	.CO(n_1027), 
	.CI(n_790), 
	.B(n_700), 
	.A(n_850));
   FAX4 g28406 (.S(n_1026), 
	.CO(n_1025), 
	.CI(n_899), 
	.B(n_840), 
	.A(n_868));
   FAX4 g28407 (.S(n_1024), 
	.CO(n_1023), 
	.CI(n_6), 
	.B(n_909), 
	.A(n_877));
   EN2X4 g28408 (.Q(n_1022), 
	.B(n_992), 
	.A(n_934));
   FAX3 g28409 (.S(n_1021), 
	.CO(n_1020), 
	.CI(n_848), 
	.B(n_664), 
	.A(n_757));
   FAX4 g28410 (.S(n_1019), 
	.CO(n_1018), 
	.CI(n_864), 
	.B(n_778), 
	.A(n_571));
   FAX4 g28411 (.S(n_1017), 
	.CO(n_1016), 
	.CI(n_898), 
	.B(n_760), 
	.A(n_687));
   FAX4 g28412 (.S(n_1015), 
	.CO(n_1014), 
	.CI(n_919), 
	.B(n_722), 
	.A(n_694));
   FAX4 g28413 (.S(n_1013), 
	.CO(n_1012), 
	.CI(n_775), 
	.B(n_876), 
	.A(n_670));
   EN3X1 g28414 (.Q(n_1011), 
	.C(n_951), 
	.B(n_934), 
	.A(n_784));
   INX4 g28415 (.Q(Z[3]), 
	.A(n_1009));
   FAX4 g28416 (.S(n_1009), 
	.CO(n_1008), 
	.CI(n_900), 
	.B(n_753), 
	.A(n_643));
   INX8 g28417 (.Q(n_1007), 
	.A(n_1006));
   FAX3 g28418 (.S(n_1006), 
	.CO(n_1005), 
	.CI(n_836), 
	.B(n_635), 
	.A(n_556));
   FAX3 g28419 (.S(n_1004), 
	.CO(n_1003), 
	.CI(n_878), 
	.B(n_459), 
	.A(n_623));
   FAX3 g28420 (.S(n_1002), 
	.CO(n_1001), 
	.CI(n_886), 
	.B(n_656), 
	.A(n_750));
   FAX4 g28421 (.S(n_1000), 
	.CO(n_999), 
	.CI(n_785), 
	.B(n_725), 
	.A(n_352));
   FAX3 g28422 (.S(n_998), 
	.CO(n_997), 
	.CI(n_852), 
	.B(n_742), 
	.A(n_520));
   FAX4 g28423 (.S(n_996), 
	.CO(n_995), 
	.CI(n_823), 
	.B(n_696), 
	.A(n_23));
   FAX4 g28424 (.S(n_994), 
	.CO(n_993), 
	.CI(n_814), 
	.B(n_748), 
	.A(n_654));
   EO2X3 g28425 (.Q(n_992), 
	.B(n_951), 
	.A(n_784));
   EN3X2 g28426 (.Q(n_991), 
	.C(n_811), 
	.B(n_692), 
	.A(n_625));
   EO2X3 g28427 (.Q(n_990), 
	.B(n_811), 
	.A(n_768));
   EO2X3 g28428 (.Q(n_989), 
	.B(n_807), 
	.A(n_771));
   EN3X2 g28429 (.Q(n_988), 
	.C(n_807), 
	.B(n_709), 
	.A(n_691));
   FAX4 g28430 (.S(n_987), 
	.CO(n_986), 
	.CI(n_754), 
	.B(n_586), 
	.A(n_649));
   FAX3 g28431 (.S(n_985), 
	.CO(n_984), 
	.CI(n_472), 
	.B(n_470), 
	.A(n_471));
   FAX4 g28432 (.S(n_983), 
	.CO(n_982), 
	.CI(n_647), 
	.B(n_648), 
	.A(n_542));
   FAX3 g28433 (.S(n_981), 
	.CO(n_980), 
	.CI(n_610), 
	.B(n_501), 
	.A(n_485));
   FAX3 g28434 (.S(n_979), 
	.CO(n_978), 
	.CI(n_461), 
	.B(n_419), 
	.A(n_460));
   FAX4 g28435 (.S(n_977), 
	.CO(n_976), 
	.CI(n_548), 
	.B(n_492), 
	.A(n_494));
   FAX3 g28436 (.S(n_975), 
	.CO(n_974), 
	.CI(n_483), 
	.B(n_424), 
	.A(n_714));
   FAX4 g28437 (.S(n_973), 
	.CO(n_972), 
	.CI(n_606), 
	.B(n_608), 
	.A(n_376));
   FAX4 g28438 (.S(n_971), 
	.CO(n_970), 
	.CI(n_776), 
	.B(n_680), 
	.A(n_679));
   FAX4 g28439 (.S(n_969), 
	.CO(n_968), 
	.CI(n_563), 
	.B(n_525), 
	.A(n_728));
   FAX4 g28440 (.S(n_967), 
	.CO(n_966), 
	.CI(n_602), 
	.B(n_726), 
	.A(n_561));
   FAX4 g28442 (.S(n_965), 
	.CO(n_964), 
	.CI(n_780), 
	.B(n_614), 
	.A(n_616));
   FAX4 g28443 (.S(n_963), 
	.CO(n_962), 
	.CI(n_701), 
	.B(n_503), 
	.A(n_663));
   FAX4 g28444 (.S(n_961), 
	.CO(n_960), 
	.CI(n_490), 
	.B(n_603), 
	.A(n_605));
   FAX3 g28445 (.S(n_959), 
	.CO(n_958), 
	.CI(n_588), 
	.B(n_734), 
	.A(n_591));
   FAX4 g28446 (.S(n_957), 
	.CO(n_956), 
	.CI(n_673), 
	.B(n_489), 
	.A(n_491));
   FAX4 g28447 (.S(n_955), 
	.CO(n_954), 
	.CI(n_580), 
	.B(n_582), 
	.A(n_584));
   FAX4 g28448 (.S(n_953), 
	.CO(n_952), 
	.CI(n_597), 
	.B(n_598), 
	.A(n_467));
   FAX4 g28449 (.S(n_951), 
	.CO(n_950), 
	.CI(n_727), 
	.B(n_517), 
	.A(n_732));
   FAX3 g28450 (.S(n_949), 
	.CO(n_948), 
	.CI(n_593), 
	.B(n_431), 
	.A(n_592));
   FAX4 g28451 (.S(n_947), 
	.CO(n_946), 
	.CI(n_569), 
	.B(n_713), 
	.A(n_358));
   INX8 g28452 (.Q(n_945), 
	.A(n_944));
   FAX3 g28453 (.S(n_944), 
	.CO(n_943), 
	.CI(n_504), 
	.B(n_374), 
	.A(n_524));
   FAX4 g28454 (.S(n_942), 
	.CO(n_941), 
	.CI(n_690), 
	.B(n_669), 
	.A(n_710));
   FAX3 g28455 (.S(n_940), 
	.CO(n_939), 
	.CI(n_533), 
	.B(n_530), 
	.A(n_697));
   FAX4 g28456 (.S(n_938), 
	.CO(n_937), 
	.CI(n_751), 
	.B(n_512), 
	.A(n_514));
   FAX4 g28457 (.S(n_936), 
	.CO(n_935), 
	.CI(n_531), 
	.B(n_535), 
	.A(n_534));
   FAX4 g28458 (.S(n_934), 
	.CO(n_933), 
	.CI(n_459), 
	.B(n_475), 
	.A(n_366));
   FAX3 g28460 (.S(n_932), 
	.CO(n_931), 
	.CI(n_510), 
	.B(n_509), 
	.A(n_507));
   FAX4 g28461 (.S(n_930), 
	.CO(n_929), 
	.CI(n_660), 
	.B(n_478), 
	.A(n_476));
   FAX3 g28462 (.S(n_928), 
	.CO(n_927), 
	.CI(n_473), 
	.B(n_526), 
	.A(n_474));
   FAX4 g28463 (.S(n_926), 
	.CO(n_925), 
	.CI(n_464), 
	.B(n_466), 
	.A(n_412));
   FAX3 g28464 (.S(n_924), 
	.CO(n_923), 
	.CI(n_540), 
	.B(n_538), 
	.A(n_537));
   FAX4 g28465 (.S(n_922), 
	.CO(n_921), 
	.CI(n_572), 
	.B(n_674), 
	.A(n_730));
   FAX3 g28467 (.S(n_920), 
	.CO(n_919), 
	.CI(n_718), 
	.B(n_370), 
	.A(n_686));
   FAX3 g28468 (.S(n_918), 
	.CO(n_917), 
	.CI(n_640), 
	.B(n_711), 
	.A(n_665));
   FAX4 g28470 (.S(n_916), 
	.CO(n_915), 
	.CI(n_611), 
	.B(n_612), 
	.A(n_415));
   FAX4 g28471 (.S(n_914), 
	.CO(n_913), 
	.CI(n_544), 
	.B(n_541), 
	.A(n_527));
   FAX3 g28472 (.S(n_912), 
	.CO(n_911), 
	.CI(n_637), 
	.B(n_368), 
	.A(n_639));
   FAX3 g28473 (.S(n_910), 
	.CO(n_909), 
	.CI(n_659), 
	.B(n_658), 
	.A(n_671));
   FAX4 g28475 (.S(n_908), 
	.CO(n_907), 
	.CI(n_559), 
	.B(n_488), 
	.A(n_486));
   FAX3 g28476 (.S(n_906), 
	.CO(n_905), 
	.CI(n_601), 
	.B(B[1]), 
	.A(n_689));
   FAX4 g28477 (.S(n_904), 
	.CO(n_903), 
	.CI(n_607), 
	.B(n_609), 
	.A(n_433));
   INX4 g28478 (.Q(Z[2]), 
	.A(n_901));
   FAX4 g28479 (.S(n_901), 
	.CO(n_900), 
	.CI(n_745), 
	.B(n_423), 
	.A(n_417));
   FAX3 g28480 (.S(n_899), 
	.CO(n_898), 
	.CI(n_468), 
	.B(n_438), 
	.A(n_573));
   FAX3 g28481 (.S(n_897), 
	.CO(n_896), 
	.CI(n_463), 
	.B(n_465), 
	.A(n_620));
   FAX3 g28482 (.S(n_895), 
	.CO(n_894), 
	.CI(n_684), 
	.B(n_583), 
	.A(n_585));
   FAX4 g28483 (.S(n_893), 
	.CO(n_892), 
	.CI(n_500), 
	.B(n_624), 
	.A(n_626));
   FAX4 g28484 (.S(n_891), 
	.CO(n_890), 
	.CI(n_733), 
	.B(n_519), 
	.A(n_576));
   FAX3 g28485 (.S(n_889), 
	.CO(n_888), 
	.CI(n_682), 
	.B(n_462), 
	.A(n_458));
   FAX4 g28486 (.S(n_887), 
	.CO(n_886), 
	.CI(n_560), 
	.B(n_421), 
	.A(n_418));
   FAX4 g28487 (.S(n_885), 
	.CO(n_884), 
	.CI(n_521), 
	.B(n_427), 
	.A(n_414));
   FAX3 g28488 (.S(n_883), 
	.CO(n_882), 
	.CI(n_545), 
	.B(n_547), 
	.A(n_543));
   FAX4 g28489 (.S(n_881), 
	.CO(n_880), 
	.CI(n_651), 
	.B(n_426), 
	.A(n_413));
   FAX3 g28490 (.S(n_879), 
	.CO(n_878), 
	.CI(n_604), 
	.B(n_22), 
	.A(n_717));
   FAX4 g28491 (.S(n_877), 
	.CO(n_876), 
	.CI(n_666), 
	.B(n_422), 
	.A(n_409));
   FAX4 g28492 (.S(n_875), 
	.CO(n_874), 
	.CI(n_642), 
	.B(n_641), 
	.A(n_442));
   FAX3 g28493 (.S(n_873), 
	.CO(n_872), 
	.CI(n_587), 
	.B(n_590), 
	.A(n_589));
   FAX3 g28494 (.S(n_871), 
	.CO(n_870), 
	.CI(n_579), 
	.B(n_578), 
	.A(n_577));
   FAX4 g28495 (.S(n_869), 
	.CO(n_868), 
	.CI(n_675), 
	.B(n_655), 
	.A(n_441));
   FAX3 g28496 (.S(n_867), 
	.CO(n_866), 
	.CI(n_532), 
	.B(n_546), 
	.A(n_539));
   FAX4 g28497 (.S(n_865), 
	.CO(n_864), 
	.CI(n_568), 
	.B(n_566), 
	.A(n_617));
   FAX3 g28498 (.S(n_863), 
	.CO(n_862), 
	.CI(n_557), 
	.B(n_554), 
	.A(n_672));
   FAX4 g28499 (.S(n_861), 
	.CO(n_860), 
	.CI(n_550), 
	.B(n_712), 
	.A(n_21));
   FAX3 g28500 (.S(n_859), 
	.CO(n_858), 
	.CI(n_564), 
	.B(n_19), 
	.A(n_721));
   FAX4 g28501 (.S(n_857), 
	.CO(n_856), 
	.CI(n_646), 
	.B(n_436), 
	.A(n_408));
   FAX4 g28503 (.S(n_855), 
	.CO(n_854), 
	.CI(n_595), 
	.B(n_522), 
	.A(n_685));
   FAX4 g28504 (.S(n_853), 
	.CO(n_852), 
	.CI(n_518), 
	.B(n_549), 
	.A(n_661));
   FAX3 g28505 (.S(n_851), 
	.CO(n_850), 
	.CI(n_716), 
	.B(n_372), 
	.A(n_699));
   FAX4 g28506 (.S(n_849), 
	.CO(n_848), 
	.CI(n_633), 
	.B(n_562), 
	.A(n_634));
   FAX4 g28507 (.S(n_847), 
	.CO(n_846), 
	.CI(n_505), 
	.B(n_506), 
	.A(n_628));
   FAX4 g28508 (.S(n_845), 
	.CO(n_844), 
	.CI(n_735), 
	.B(n_515), 
	.A(n_378));
   FAX4 g28509 (.S(n_843), 
	.CO(n_842), 
	.CI(n_691), 
	.B(n_599), 
	.A(n_715));
   FAX3 g28510 (.S(n_841), 
	.CO(n_840), 
	.CI(n_574), 
	.B(n_411), 
	.A(n_516));
   FAX4 g28511 (.S(n_839), 
	.CO(n_838), 
	.CI(n_487), 
	.B(n_719), 
	.A(n_362));
   FAX4 g28512 (.S(n_837), 
	.CO(n_836), 
	.CI(n_498), 
	.B(n_706), 
	.A(n_497));
   INX8 g28513 (.Q(n_835), 
	.A(n_834));
   FAX3 g28514 (.S(n_834), 
	.CO(n_833), 
	.CI(n_703), 
	.B(n_354), 
	.A(n_484));
   FAX3 g28515 (.S(n_832), 
	.CO(n_831), 
	.CI(n_683), 
	.B(n_18), 
	.A(n_705));
   FAX3 g28516 (.S(n_830), 
	.CO(n_829), 
	.CI(n_558), 
	.B(n_618), 
	.A(n_596));
   FAX4 g28517 (.S(n_828), 
	.CO(n_827), 
	.CI(n_482), 
	.B(n_481), 
	.A(n_630));
   FAX4 g28518 (.S(n_826), 
	.CO(n_825), 
	.CI(n_681), 
	.B(n_678), 
	.A(n_551));
   FAX3 g28519 (.S(n_824), 
	.CO(n_823), 
	.CI(n_496), 
	.B(n_650), 
	.A(n_645));
   FAX3 g28520 (.S(n_822), 
	.CO(n_821), 
	.CI(n_567), 
	.B(n_570), 
	.A(n_738));
   FAX4 g28521 (.S(n_820), 
	.CO(n_819), 
	.CI(n_638), 
	.B(n_704), 
	.A(n_25));
   FAX4 g28522 (.S(n_818), 
	.CO(n_817), 
	.CI(n_631), 
	.B(n_668), 
	.A(n_432));
   FAX4 g28523 (.S(n_816), 
	.CO(n_815), 
	.CI(n_552), 
	.B(n_429), 
	.A(n_416));
   FAX3 g28524 (.S(n_814), 
	.CO(n_813), 
	.CI(n_657), 
	.B(n_410), 
	.A(n_440));
   EN3X2 g28525 (.Q(n_812), 
	.C(n_575), 
	.B(n_581), 
	.A(n_382));
   EN3X1 g28527 (.Q(n_811), 
	.C(n_621), 
	.B(n_720), 
	.A(n_622));
   EN2X4 g28528 (.Q(n_810), 
	.B(n_765), 
	.A(n_720));
   EN3X2 g28529 (.Q(n_809), 
	.C(n_652), 
	.B(n_536), 
	.A(n_737));
   EN3X2 g28530 (.Q(n_808), 
	.C(n_513), 
	.B(n_511), 
	.A(n_731));
   EN3X1 g28531 (.Q(n_807), 
	.C(n_667), 
	.B(n_502), 
	.A(n_739));
   EN2X4 g28532 (.Q(n_806), 
	.B(n_770), 
	.A(n_644));
   EN3X1 g28533 (.Q(n_805), 
	.C(n_615), 
	.B(n_613), 
	.A(n_600));
   EN3X1 g28534 (.Q(n_804), 
	.C(n_495), 
	.B(n_508), 
	.A(n_688));
   EN3X2 g28535 (.Q(n_803), 
	.C(n_479), 
	.B(n_480), 
	.A(n_477));
   EN2X4 g28536 (.Q(n_802), 
	.B(n_763), 
	.A(n_667));
   EO2X3 g28537 (.Q(n_801), 
	.B(n_761), 
	.A(n_511));
   EO2X3 g28538 (.Q(n_800), 
	.B(n_762), 
	.A(n_652));
   EN3X1 g28539 (.Q(n_799), 
	.C(n_644), 
	.B(n_565), 
	.A(n_724));
   EN2X4 g28540 (.Q(n_798), 
	.B(n_767), 
	.A(n_495));
   EO2X3 g28541 (.Q(n_797), 
	.B(n_766), 
	.A(n_477));
   EN2X4 g28542 (.Q(n_796), 
	.B(n_764), 
	.A(n_613));
   EN3X2 g28543 (.Q(n_795), 
	.C(n_746), 
	.B(n_619), 
	.A(n_662));
   EN3X2 g28544 (.Q(n_794), 
	.C(n_553), 
	.B(n_743), 
	.A(n_555));
   EN3X2 g28545 (.Q(n_793), 
	.C(n_740), 
	.B(n_627), 
	.A(n_469));
   EN2X4 g28546 (.Q(n_792), 
	.B(n_772), 
	.A(n_352));
   EN2X4 g28551 (.Q(n_791), 
	.B(n_774), 
	.A(n_499));
   EN3X1 g28553 (.Q(n_790), 
	.C(n_707), 
	.B(n_736), 
	.A(n_364));
   EN2X4 g28554 (.Q(n_789), 
	.B(n_779), 
	.A(n_698));
   EN3X2 g28555 (.Q(n_788), 
	.C(n_632), 
	.B(n_381), 
	.A(n_653));
   EN3X1 g28556 (.Q(n_787), 
	.C(n_523), 
	.B(n_499), 
	.A(n_20));
   EN3X2 g28557 (.Q(n_786), 
	.C(n_528), 
	.B(n_493), 
	.A(n_356));
   EN3X2 g28558 (.Q(n_785), 
	.C(n_708), 
	.B(n_364), 
	.A(n_736));
   EN3X2 g28559 (.Q(n_784), 
	.C(n_723), 
	.B(n_698), 
	.A(n_24));
   EN2X4 g28560 (.Q(n_783), 
	.B(n_493), 
	.A(n_356));
   EN2X4 g28561 (.Q(n_782), 
	.B(n_662), 
	.A(n_619));
   EN2X4 g28562 (.Q(n_781), 
	.B(n_632), 
	.A(n_381));
   EN2X4 g28563 (.Q(n_780), 
	.B(n_629), 
	.A(n_447));
   EN2X4 g28564 (.Q(n_779), 
	.B(n_723), 
	.A(n_24));
   EN2X4 g28565 (.Q(n_778), 
	.B(n_594), 
	.A(n_451));
   EO2X3 g28566 (.Q(n_777), 
	.B(n_553), 
	.A(n_555));
   EN2X4 g28567 (.Q(n_776), 
	.B(n_529), 
	.A(n_457));
   EN2X4 g28568 (.Q(n_775), 
	.B(n_636), 
	.A(n_456));
   EO2X3 g28569 (.Q(n_774), 
	.B(n_523), 
	.A(n_20));
   EN2X4 g28570 (.Q(n_773), 
	.B(n_627), 
	.A(n_469));
   EO2X3 g28571 (.Q(n_772), 
	.B(n_729), 
	.A(n_360));
   EO2X3 g28572 (.Q(n_771), 
	.B(n_691), 
	.A(n_709));
   EO2X3 g28573 (.Q(n_770), 
	.B(n_565), 
	.A(n_724));
   EO2X3 g28574 (.Q(n_769), 
	.B(n_581), 
	.A(n_382));
   EO2X3 g28575 (.Q(n_768), 
	.B(n_692), 
	.A(n_625));
   EO2X3 g28576 (.Q(n_767), 
	.B(n_508), 
	.A(n_688));
   EO2X3 g28577 (.Q(n_766), 
	.B(n_479), 
	.A(n_480));
   EO2X3 g28578 (.Q(n_765), 
	.B(n_621), 
	.A(n_622));
   EO2X3 g28579 (.Q(n_764), 
	.B(n_615), 
	.A(n_600));
   EO2X3 g28580 (.Q(n_763), 
	.B(n_502), 
	.A(n_739));
   EO2X3 g28581 (.Q(n_762), 
	.B(n_536), 
	.A(n_737));
   EO2X3 g28582 (.Q(n_761), 
	.B(n_513), 
	.A(n_731));
   OR2X4 g28583 (.Q(n_760), 
	.B(n_529), 
	.A(n_457));
   OR2X4 g28584 (.Q(n_759), 
	.B(n_636), 
	.A(n_456));
   OR2X4 g28585 (.Q(n_758), 
	.B(n_594), 
	.A(n_451));
   OR2X4 g28586 (.Q(n_757), 
	.B(n_629), 
	.A(n_447));
   AN21X4 g28587 (.Q(Z[1]), 
	.C(n_744), 
	.B(n_435), 
	.A(n_340));
   EN2X4 g28588 (.Q(n_755), 
	.B(n_434), 
	.A(n_453));
   EN2X4 g28589 (.Q(n_754), 
	.B(n_437), 
	.A(n_452));
   EN2X4 g28590 (.Q(n_753), 
	.B(n_439), 
	.A(n_455));
   EN2X4 g28591 (.Q(n_752), 
	.B(n_430), 
	.A(n_454));
   EN2X4 g28592 (.Q(n_751), 
	.B(n_425), 
	.A(n_448));
   EN2X4 g28593 (.Q(n_750), 
	.B(n_428), 
	.A(n_449));
   EN2X4 g28594 (.Q(n_749), 
	.B(n_420), 
	.A(n_450));
   OR2X4 g28595 (.Q(n_748), 
	.B(n_437), 
	.A(n_452));
   OR2X4 g28596 (.Q(n_747), 
	.B(n_439), 
	.A(n_455));
   NO2X4 g28597 (.Q(n_746), 
	.B(n_434), 
	.A(n_453));
   INX8 g28598 (.Q(n_745), 
	.A(n_744));
   NO2X4 g28599 (.Q(n_744), 
	.B(n_435), 
	.A(n_340));
   NO2X4 g28600 (.Q(n_743), 
	.B(n_430), 
	.A(n_454));
   OR2X4 g28601 (.Q(n_742), 
	.B(n_425), 
	.A(n_448));
   OR2X4 g28602 (.Q(n_741), 
	.B(n_428), 
	.A(n_449));
   NO2X4 g28603 (.Q(n_740), 
	.B(n_420), 
	.A(n_450));
   ON21X4 g28604 (.Q(n_739), 
	.C(B[9]), 
	.B(n_385), 
	.A(n_88));
   AN21X2  g28605 (.Q(n_738), 
	.C(n_17), 
	.B(n_394), 
	.A(n_186));
   AN21X2  g28606 (.Q(n_737), 
	.C(n_15), 
	.B(n_395), 
	.A(n_100));
   ON21X4 g28607 (.Q(n_736), 
	.C(B[21]), 
	.B(n_387), 
	.A(n_174));
   ON21X4 g28608 (.Q(n_735), 
	.C(B[19]), 
	.B(n_404), 
	.A(n_66));
   ON21X4 g28609 (.Q(n_734), 
	.C(B[5]), 
	.B(n_390), 
	.A(n_96));
   AN21X2  g28610 (.Q(n_733), 
	.C(n_16), 
	.B(n_388), 
	.A(n_182));
   ON21X4 g28611 (.Q(n_732), 
	.C(B[17]), 
	.B(n_406), 
	.A(n_119));
   AN21X2  g28612 (.Q(n_731), 
	.C(n_14), 
	.B(n_392), 
	.A(n_305));
   AN21X2  g28613 (.Q(n_730), 
	.C(n_13), 
	.B(n_401), 
	.A(n_266));
   ON21X4 g28614 (.Q(n_729), 
	.C(B[23]), 
	.B(n_397), 
	.A(n_2));
   AN22X2 g28615 (.Q(n_728), 
	.D(n_2), 
	.C(n_355), 
	.B(n_397), 
	.A(n_27));
   AO22X4 g28616 (.Q(n_727), 
	.D(n_2), 
	.C(n_379), 
	.B(n_397), 
	.A(n_371));
   AN22X2 g28617 (.Q(n_726), 
	.D(n_2), 
	.C(n_28), 
	.B(n_397), 
	.A(n_375));
   AN22X2 g28618 (.Q(n_725), 
	.D(B[23]), 
	.C(n_2), 
	.B(n_397), 
	.A(n_361));
   AO22X4 g28619 (.Q(n_724), 
	.D(n_2), 
	.C(n_26), 
	.B(n_397), 
	.A(n_363));
   AN22X2 g28620 (.Q(n_723), 
	.D(n_371), 
	.C(n_2), 
	.B(n_397), 
	.A(n_367));
   AO22X4 g28621 (.Q(n_722), 
	.D(n_2), 
	.C(n_365), 
	.B(n_397), 
	.A(n_373));
   AN22X2 g28622 (.Q(n_721), 
	.D(n_357), 
	.C(n_2), 
	.B(n_397), 
	.A(n_33));
   AN22X2 g28623 (.Q(n_720), 
	.D(n_2), 
	.C(n_363), 
	.B(n_397), 
	.A(n_369));
   AO22X4 g28624 (.Q(n_719), 
	.D(n_2), 
	.C(n_31), 
	.B(n_397), 
	.A(n_26));
   AO22X4 g28625 (.Q(n_718), 
	.D(n_2), 
	.C(n_373), 
	.B(n_397), 
	.A(n_379));
   AN22X2 g28626 (.Q(n_717), 
	.D(n_367), 
	.C(n_2), 
	.B(n_397), 
	.A(n_32));
   AO22X4 g28627 (.Q(n_716), 
	.D(n_2), 
	.C(n_353), 
	.B(n_397), 
	.A(n_365));
   AN22X2 g28628 (.Q(n_715), 
	.D(n_2), 
	.C(n_33), 
	.B(n_397), 
	.A(n_30));
   AN22X2 g28629 (.Q(n_714), 
	.D(n_2), 
	.C(n_27), 
	.B(n_397), 
	.A(n_380));
   AO22X4 g28630 (.Q(n_713), 
	.D(n_2), 
	.C(n_369), 
	.B(n_397), 
	.A(n_377));
   AN22X2 g28631 (.Q(n_712), 
	.D(n_377), 
	.C(n_2), 
	.B(n_397), 
	.A(n_359));
   AN22X2 g28632 (.Q(n_711), 
	.D(n_29), 
	.C(n_2), 
	.B(n_397), 
	.A(n_357));
   AN22X2 g28633 (.Q(n_710), 
	.D(n_2), 
	.C(n_32), 
	.B(n_397), 
	.A(n_29));
   AO22X4 g28634 (.Q(n_709), 
	.D(n_2), 
	.C(n_30), 
	.B(n_397), 
	.A(n_383));
   INX4 g28635 (.Q(n_708), 
	.A(n_707));
   AN22X2 g28636 (.Q(n_707), 
	.D(n_361), 
	.C(n_2), 
	.B(n_397), 
	.A(n_353));
   AN22X2 g28637 (.Q(n_706), 
	.D(n_2), 
	.C(n_359), 
	.B(n_397), 
	.A(n_28));
   AN22X2 g28638 (.Q(n_705), 
	.D(n_383), 
	.C(n_2), 
	.B(n_397), 
	.A(n_31));
   AN22X2 g28639 (.Q(n_704), 
	.D(n_2), 
	.C(n_375), 
	.B(n_397), 
	.A(n_355));
   ON22X4 g28640 (.Q(n_703), 
	.D(n_305), 
	.C(n_14), 
	.B(n_392), 
	.A(n_106));
   INX8 g28641 (.Q(n_702), 
	.A(n_701));
   AN22X2 g28642 (.Q(n_701), 
	.D(n_88), 
	.C(B[9]), 
	.B(n_385), 
	.A(n_40));
   INX8 g28643 (.Q(n_700), 
	.A(n_699));
   AN22X2 g28644 (.Q(n_699), 
	.D(B[21]), 
	.C(n_174), 
	.B(n_387), 
	.A(n_178));
   AN22X2 g28645 (.Q(n_698), 
	.D(n_119), 
	.C(B[17]), 
	.B(n_406), 
	.A(n_246));
   AN22X2 g28646 (.Q(n_697), 
	.D(B[5]), 
	.C(n_96), 
	.B(n_390), 
	.A(n_258));
   INX8 g28647 (.Q(n_696), 
	.A(n_695));
   ON22X4 g28648 (.Q(n_695), 
	.D(n_266), 
	.C(n_13), 
	.B(n_401), 
	.A(n_76));
   INX8 g28649 (.Q(n_694), 
	.A(n_693));
   AN22X2 g28650 (.Q(n_693), 
	.D(n_66), 
	.C(B[19]), 
	.B(n_404), 
	.A(n_212));
   OA22X4 g28651 (.Q(n_692), 
	.D(n_100), 
	.C(n_15), 
	.B(n_395), 
	.A(n_291));
   OA22X4 g28652 (.Q(n_691), 
	.D(n_186), 
	.C(n_17), 
	.B(n_394), 
	.A(n_47));
   AN22X2 g28653 (.Q(n_690), 
	.D(B[15]), 
	.C(n_183), 
	.B(n_389), 
	.A(n_77));
   AN22X2 g28654 (.Q(n_689), 
	.D(n_147), 
	.C(n_267), 
	.B(n_402), 
	.A(n_152));
   ON22X4 g28655 (.Q(n_688), 
	.D(n_65), 
	.C(n_158), 
	.B(n_403), 
	.A(n_143));
   AN22X2 g28656 (.Q(n_687), 
	.D(n_96), 
	.C(n_167), 
	.B(n_390), 
	.A(n_99));
   ON22X4 g28657 (.Q(n_686), 
	.D(n_173), 
	.C(n_160), 
	.B(n_386), 
	.A(n_286));
   AN22X2 g28658 (.Q(n_685), 
	.D(n_119), 
	.C(n_130), 
	.B(n_406), 
	.A(n_109));
   AN22X2 g28659 (.Q(n_684), 
	.D(n_138), 
	.C(n_101), 
	.B(n_396), 
	.A(n_256));
   AN22X2 g28660 (.Q(n_683), 
	.D(n_63), 
	.C(n_119), 
	.B(n_406), 
	.A(n_104));
   AN22X2 g28661 (.Q(n_682), 
	.D(n_191), 
	.C(n_267), 
	.B(n_402), 
	.A(n_131));
   AN22X2 g28662 (.Q(n_681), 
	.D(n_216), 
	.C(n_96), 
	.B(n_390), 
	.A(n_288));
   AN22X2 g28663 (.Q(n_680), 
	.D(n_96), 
	.C(n_99), 
	.B(n_390), 
	.A(n_151));
   OA22X4 g28664 (.Q(n_679), 
	.D(n_186), 
	.C(n_232), 
	.B(n_394), 
	.A(n_322));
   AN22X2 g28665 (.Q(n_678), 
	.D(n_88), 
	.C(n_284), 
	.B(n_385), 
	.A(n_210));
   INX8 g28666 (.Q(n_677), 
	.A(n_676));
   ON22X4 g28667 (.Q(n_676), 
	.D(n_305), 
	.C(n_106), 
	.B(n_392), 
	.A(n_289));
   AN22X2 g28668 (.Q(n_675), 
	.D(n_151), 
	.C(n_96), 
	.B(n_390), 
	.A(n_224));
   AN22X2 g28669 (.Q(n_674), 
	.D(n_77), 
	.C(n_183), 
	.B(n_389), 
	.A(n_145));
   AN22X2 g28670 (.Q(n_673), 
	.D(n_85), 
	.C(n_88), 
	.B(n_385), 
	.A(n_122));
   AN22X2 g28671 (.Q(n_672), 
	.D(n_43), 
	.C(n_183), 
	.B(n_389), 
	.A(n_222));
   AN22X2 g28672 (.Q(n_671), 
	.D(n_244), 
	.C(n_96), 
	.B(n_390), 
	.A(n_206));
   AN22X2 g28673 (.Q(n_670), 
	.D(n_96), 
	.C(n_224), 
	.B(n_390), 
	.A(n_176));
   AN22X2 g28674 (.Q(n_669), 
	.D(n_144), 
	.C(n_174), 
	.B(n_387), 
	.A(n_153));
   AN22X2 g28675 (.Q(n_668), 
	.D(n_88), 
	.C(n_41), 
	.B(n_385), 
	.A(n_328));
   ON22X4 g28676 (.Q(n_667), 
	.D(n_182), 
	.C(n_282), 
	.B(n_388), 
	.A(n_169));
   AN22X2 g28677 (.Q(n_666), 
	.D(n_101), 
	.C(n_93), 
	.B(n_396), 
	.A(n_255));
   AN22X2 g28678 (.Q(n_665), 
	.D(n_153), 
	.C(n_174), 
	.B(n_387), 
	.A(n_141));
   AN22X2 g28679 (.Q(n_664), 
	.D(n_152), 
	.C(n_267), 
	.B(n_402), 
	.A(n_215));
   ON22X4 g28680 (.Q(n_663), 
	.D(n_173), 
	.C(n_277), 
	.B(n_386), 
	.A(n_56));
   ON22X4 g28681 (.Q(n_662), 
	.D(n_305), 
	.C(n_263), 
	.B(n_392), 
	.A(n_39));
   AN22X2 g28682 (.Q(n_661), 
	.D(n_119), 
	.C(n_109), 
	.B(n_406), 
	.A(n_319));
   AN22X2 g28683 (.Q(n_660), 
	.D(n_51), 
	.C(n_96), 
	.B(n_390), 
	.A(n_167));
   OA22X4 g28684 (.Q(n_659), 
	.D(n_305), 
	.C(n_39), 
	.B(n_392), 
	.A(n_195));
   AN22X2 g28685 (.Q(n_658), 
	.D(n_101), 
	.C(n_255), 
	.B(n_396), 
	.A(n_320));
   OA22X4 g28686 (.Q(n_657), 
	.D(n_305), 
	.C(n_195), 
	.B(n_392), 
	.A(n_187));
   AN22X2 g28687 (.Q(n_656), 
	.D(n_53), 
	.C(n_267), 
	.B(n_402), 
	.A(n_181));
   AN22X2 g28688 (.Q(n_655), 
	.D(n_88), 
	.C(n_81), 
	.B(n_385), 
	.A(n_41));
   AN22X2 g28689 (.Q(n_654), 
	.D(n_96), 
	.C(n_206), 
	.B(n_390), 
	.A(n_253));
   AO22X4 g28690 (.Q(n_653), 
	.D(n_101), 
	.C(n_256), 
	.B(n_396), 
	.A(n_225));
   AN22X2 g28691 (.Q(n_652), 
	.D(n_267), 
	.C(n_73), 
	.B(n_402), 
	.A(n_290));
   AN22X2 g28692 (.Q(n_651), 
	.D(n_247), 
	.C(n_304), 
	.B(n_391), 
	.A(n_155));
   AN22X2 g28693 (.Q(n_650), 
	.D(n_141), 
	.C(n_174), 
	.B(n_387), 
	.A(n_184));
   AN22X2 g28694 (.Q(n_649), 
	.D(n_96), 
	.C(n_253), 
	.B(n_390), 
	.A(n_324));
   AN22X2 g28695 (.Q(n_648), 
	.D(n_183), 
	.C(n_128), 
	.B(n_389), 
	.A(n_211));
   AN22X2 g28696 (.Q(n_647), 
	.D(n_35), 
	.C(n_88), 
	.B(n_385), 
	.A(n_261));
   AN22X2 g28697 (.Q(n_646), 
	.D(n_304), 
	.C(n_146), 
	.B(n_391), 
	.A(n_162));
   AN22X2 g28698 (.Q(n_645), 
	.D(n_145), 
	.C(n_183), 
	.B(n_389), 
	.A(n_189));
   ON22X4 g28699 (.Q(n_644), 
	.D(n_182), 
	.C(n_59), 
	.B(n_388), 
	.A(n_124));
   AN22X2 g28700 (.Q(n_643), 
	.D(n_304), 
	.C(n_162), 
	.B(n_391), 
	.A(n_326));
   AN22X2 g28701 (.Q(n_642), 
	.D(n_132), 
	.C(n_66), 
	.B(n_404), 
	.A(n_117));
   AN22X2 g28702 (.Q(n_641), 
	.D(n_174), 
	.C(n_285), 
	.B(n_387), 
	.A(n_237));
   AN22X2 g28703 (.Q(n_640), 
	.D(n_273), 
	.C(n_119), 
	.B(n_406), 
	.A(n_243));
   ON22X4 g28704 (.Q(n_639), 
	.D(n_118), 
	.C(n_202), 
	.B(n_405), 
	.A(n_136));
   AN22X2 g28705 (.Q(n_638), 
	.D(n_259), 
	.C(n_3), 
	.B(n_393), 
	.A(n_270));
   ON22X4 g28706 (.Q(n_637), 
	.D(n_186), 
	.C(n_45), 
	.B(n_394), 
	.A(n_114));
   OA22X4 g28707 (.Q(n_636), 
	.D(n_305), 
	.C(n_46), 
	.B(n_392), 
	.A(n_263));
   AN22X2 g28708 (.Q(n_635), 
	.D(n_140), 
	.C(n_119), 
	.B(n_406), 
	.A(n_257));
   AN22X2 g28709 (.Q(n_634), 
	.D(n_174), 
	.C(n_237), 
	.B(n_387), 
	.A(n_203));
   AN22X2 g28710 (.Q(n_633), 
	.D(n_261), 
	.C(n_88), 
	.B(n_385), 
	.A(n_200));
   ON22X4 g28711 (.Q(n_632), 
	.D(n_305), 
	.C(n_289), 
	.B(n_392), 
	.A(n_207));
   AN22X2 g28712 (.Q(n_631), 
	.D(n_101), 
	.C(n_86), 
	.B(n_396), 
	.A(n_93));
   AN22X2 g28713 (.Q(n_630), 
	.D(n_88), 
	.C(n_219), 
	.B(n_385), 
	.A(n_61));
   OA22X4 g28714 (.Q(n_629), 
	.D(n_305), 
	.C(n_207), 
	.B(n_392), 
	.A(n_209));
   AN22X2 g28715 (.Q(n_628), 
	.D(n_88), 
	.C(n_92), 
	.B(n_385), 
	.A(n_85));
   ON22X4 g28716 (.Q(n_627), 
	.D(n_186), 
	.C(n_251), 
	.B(n_394), 
	.A(n_179));
   AN22X2 g28717 (.Q(n_626), 
	.D(n_119), 
	.C(n_90), 
	.B(n_406), 
	.A(n_214));
   AN22X2 g28718 (.Q(n_625), 
	.D(n_66), 
	.C(n_97), 
	.B(n_404), 
	.A(n_201));
   AN22X2 g28719 (.Q(n_624), 
	.D(n_183), 
	.C(n_211), 
	.B(n_389), 
	.A(n_205));
   AN22X2 g28720 (.Q(n_623), 
	.D(n_120), 
	.C(n_174), 
	.B(n_387), 
	.A(n_172));
   AN22X2 g28721 (.Q(n_622), 
	.D(n_174), 
	.C(n_111), 
	.B(n_387), 
	.A(n_236));
   AN22X2 g28722 (.Q(n_621), 
	.D(n_267), 
	.C(n_290), 
	.B(n_402), 
	.A(n_208));
   AN22X2 g28723 (.Q(n_620), 
	.D(n_262), 
	.C(n_66), 
	.B(n_404), 
	.A(n_132));
   AO22X4 g28724 (.Q(n_619), 
	.D(n_96), 
	.C(n_176), 
	.B(n_390), 
	.A(n_244));
   AN22X2 g28725 (.Q(n_618), 
	.D(n_78), 
	.C(n_267), 
	.B(n_402), 
	.A(n_147));
   AN22X2 g28726 (.Q(n_617), 
	.D(n_119), 
	.C(n_241), 
	.B(n_406), 
	.A(n_220));
   AN22X2 g28727 (.Q(n_616), 
	.D(n_267), 
	.C(n_215), 
	.B(n_402), 
	.A(n_67));
   ON22X4 g28728 (.Q(n_615), 
	.D(n_186), 
	.C(n_114), 
	.B(n_394), 
	.A(n_196));
   AN22X2 g28729 (.Q(n_614), 
	.D(n_3), 
	.C(n_234), 
	.B(n_393), 
	.A(n_197));
   AO22X4 g28730 (.Q(n_613), 
	.D(n_66), 
	.C(n_201), 
	.B(n_404), 
	.A(n_107));
   AN22X2 g28731 (.Q(n_612), 
	.D(n_161), 
	.C(n_101), 
	.B(n_396), 
	.A(n_135));
   OA22X4 g28732 (.Q(n_611), 
	.D(n_305), 
	.C(n_209), 
	.B(n_392), 
	.A(n_194));
   AN22X2 g28733 (.Q(n_610), 
	.D(n_80), 
	.C(n_96), 
	.B(n_390), 
	.A(n_250));
   AN22X2 g28734 (.Q(n_609), 
	.D(n_174), 
	.C(n_203), 
	.B(n_387), 
	.A(n_127));
   ON22X4 g28735 (.Q(n_608), 
	.D(n_87), 
	.C(n_265), 
	.B(n_384), 
	.A(n_192));
   AN22X2 g28736 (.Q(n_607), 
	.D(n_264), 
	.C(n_66), 
	.B(n_404), 
	.A(n_193));
   ON22X4 g28737 (.Q(n_606), 
	.D(n_182), 
	.C(n_124), 
	.B(n_388), 
	.A(n_44));
   AN22X2 g28738 (.Q(n_605), 
	.D(n_3), 
	.C(n_197), 
	.B(n_393), 
	.A(n_190));
   AN22X2 g28739 (.Q(n_604), 
	.D(n_223), 
	.C(n_66), 
	.B(n_404), 
	.A(n_149));
   AN22X2 g28740 (.Q(n_603), 
	.D(n_267), 
	.C(n_67), 
	.B(n_402), 
	.A(n_165));
   AN22X2 g28741 (.Q(n_602), 
	.D(n_274), 
	.C(n_3), 
	.B(n_393), 
	.A(n_259));
   AN22X2 g28742 (.Q(n_601), 
	.D(n_276), 
	.C(n_96), 
	.B(n_390), 
	.A(n_171));
   ON22X4 g28743 (.Q(n_600), 
	.D(n_118), 
	.C(n_136), 
	.B(n_405), 
	.A(n_37));
   AN22X2 g28744 (.Q(n_599), 
	.D(n_184), 
	.C(n_174), 
	.B(n_387), 
	.A(n_94));
   AN22X2 g28745 (.Q(n_598), 
	.D(n_183), 
	.C(n_205), 
	.B(n_389), 
	.A(n_175));
   AN22X2 g28746 (.Q(n_597), 
	.D(n_200), 
	.C(n_88), 
	.B(n_385), 
	.A(n_91));
   AN22X2 g28747 (.Q(n_596), 
	.D(n_115), 
	.C(n_183), 
	.B(n_389), 
	.A(n_55));
   AN22X2 g28748 (.Q(n_595), 
	.D(n_260), 
	.C(n_304), 
	.B(n_391), 
	.A(n_272));
   OA22X4 g28749 (.Q(n_594), 
	.D(n_305), 
	.C(n_194), 
	.B(n_392), 
	.A(n_188));
   AN22X2 g28750 (.Q(n_593), 
	.D(n_89), 
	.C(n_96), 
	.B(n_390), 
	.A(n_216));
   AN22X2 g28751 (.Q(n_592), 
	.D(n_190), 
	.C(n_3), 
	.B(n_393), 
	.A(n_168));
   ON22X4 g28752 (.Q(n_591), 
	.D(n_100), 
	.C(n_291), 
	.B(n_395), 
	.A(n_34));
   AN22X2 g28753 (.Q(n_590), 
	.D(n_174), 
	.C(n_127), 
	.B(n_387), 
	.A(n_323));
   AN22X2 g28754 (.Q(n_589), 
	.D(n_66), 
	.C(n_193), 
	.B(n_404), 
	.A(n_113));
   ON22X4 g28755 (.Q(n_588), 
	.D(n_186), 
	.C(n_196), 
	.B(n_394), 
	.A(n_98));
   AN22X2 g28756 (.Q(n_587), 
	.D(n_91), 
	.C(n_88), 
	.B(n_385), 
	.A(n_284));
   AN21X4 g28757 (.Q(n_586), 
	.C(n_407), 
	.B(n_391), 
	.A(n_146));
   AN22X2 g28758 (.Q(n_585), 
	.D(n_55), 
	.C(n_183), 
	.B(n_389), 
	.A(n_128));
   AO22X4 g28759 (.Q(n_584), 
	.D(n_174), 
	.C(n_236), 
	.B(n_387), 
	.A(n_185));
   AN22X2 g28760 (.Q(n_583), 
	.D(n_119), 
	.C(n_133), 
	.B(n_406), 
	.A(n_279));
   AO22X4 g28761 (.Q(n_582), 
	.D(n_66), 
	.C(n_107), 
	.B(n_404), 
	.A(n_110));
   ON22X4 g28762 (.Q(n_581), 
	.D(n_65), 
	.C(n_48), 
	.B(n_403), 
	.A(n_159));
   AO22X4 g28763 (.Q(n_580), 
	.D(n_267), 
	.C(n_208), 
	.B(n_402), 
	.A(n_38));
   AN22X2 g28764 (.Q(n_579), 
	.D(n_135), 
	.C(n_101), 
	.B(n_396), 
	.A(n_50));
   AN22X2 g28765 (.Q(n_578), 
	.D(n_52), 
	.C(n_119), 
	.B(n_406), 
	.A(n_241));
   AN22X2 g28766 (.Q(n_577), 
	.D(n_175), 
	.C(n_183), 
	.B(n_389), 
	.A(n_157));
   AN22X2 g28767 (.Q(n_576), 
	.D(n_119), 
	.C(n_246), 
	.B(n_406), 
	.A(n_62));
   AO22X4 g28768 (.Q(n_575), 
	.D(n_183), 
	.C(n_189), 
	.B(n_389), 
	.A(n_71));
   OA22X4 g28769 (.Q(n_574), 
	.D(n_305), 
	.C(n_134), 
	.B(n_392), 
	.A(n_46));
   AN22X2 g28770 (.Q(n_573), 
	.D(n_88), 
	.C(n_64), 
	.B(n_385), 
	.A(n_81));
   AN22X2 g28771 (.Q(n_572), 
	.D(n_102), 
	.C(n_66), 
	.B(n_404), 
	.A(n_83));
   AN22X2 g28772 (.Q(n_571), 
	.D(n_267), 
	.C(n_165), 
	.B(n_402), 
	.A(n_156));
   AN22X2 g28773 (.Q(n_570), 
	.D(n_242), 
	.C(n_119), 
	.B(n_406), 
	.A(n_170));
   ON22X4 g28774 (.Q(n_569), 
	.D(n_87), 
	.C(n_192), 
	.B(n_384), 
	.A(n_240));
   OA22X4 g28775 (.Q(n_568), 
	.D(n_305), 
	.C(n_188), 
	.B(n_392), 
	.A(n_108));
   OA22X4 g28776 (.Q(n_567), 
	.D(n_266), 
	.C(n_76), 
	.B(n_401), 
	.A(n_148));
   AN22X2 g28777 (.Q(n_566), 
	.D(n_157), 
	.C(n_183), 
	.B(n_389), 
	.A(n_150));
   ON22X4 g28778 (.Q(n_565), 
	.D(n_173), 
	.C(n_56), 
	.B(n_386), 
	.A(n_112));
   AN22X2 g28779 (.Q(n_564), 
	.D(n_243), 
	.C(n_119), 
	.B(n_406), 
	.A(n_242));
   AN22X2 g28780 (.Q(n_563), 
	.D(n_171), 
	.C(n_96), 
	.B(n_390), 
	.A(n_271));
   AN22X2 g28781 (.Q(n_562), 
	.D(n_66), 
	.C(n_117), 
	.B(n_404), 
	.A(n_264));
   AN22X2 g28782 (.Q(n_561), 
	.D(n_174), 
	.C(n_79), 
	.B(n_387), 
	.A(n_252));
   AN22X2 g28783 (.Q(n_560), 
	.D(n_235), 
	.C(n_304), 
	.B(n_391), 
	.A(n_72));
   AN22X2 g28784 (.Q(n_559), 
	.D(n_155), 
	.C(n_304), 
	.B(n_391), 
	.A(n_235));
   AO22X4 g28785 (.Q(n_558), 
	.D(n_96), 
	.C(n_58), 
	.B(n_390), 
	.A(n_276));
   INX8 g28786 (.Q(n_557), 
	.A(n_556));
   ON22X4 g28787 (.Q(n_556), 
	.D(n_100), 
	.C(n_34), 
	.B(n_395), 
	.A(n_142));
   AO22X4 g28788 (.Q(n_555), 
	.D(n_267), 
	.C(n_156), 
	.B(n_402), 
	.A(n_217));
   AN22X2 g28789 (.Q(n_554), 
	.D(n_36), 
	.C(n_119), 
	.B(n_406), 
	.A(n_140));
   AO22X4 g28790 (.Q(n_553), 
	.D(n_3), 
	.C(n_168), 
	.B(n_393), 
	.A(n_126));
   AN22X2 g28791 (.Q(n_552), 
	.D(n_50), 
	.C(n_101), 
	.B(n_396), 
	.A(n_198));
   AN22X2 g28792 (.Q(n_551), 
	.D(n_66), 
	.C(n_113), 
	.B(n_404), 
	.A(n_123));
   AN22X2 g28793 (.Q(n_550), 
	.D(n_38), 
	.C(n_267), 
	.B(n_402), 
	.A(n_218));
   AN22X2 g28794 (.Q(n_549), 
	.D(n_183), 
	.C(n_70), 
	.B(n_389), 
	.A(n_228));
   AN22X2 g28795 (.Q(n_548), 
	.D(n_69), 
	.C(n_96), 
	.B(n_390), 
	.A(n_80));
   AN22X2 g28796 (.Q(n_547), 
	.D(n_220), 
	.C(n_119), 
	.B(n_406), 
	.A(n_130));
   AN22X2 g28797 (.Q(n_546), 
	.D(n_94), 
	.C(n_174), 
	.B(n_387), 
	.A(n_238));
   AN22X2 g28798 (.Q(n_545), 
	.D(n_198), 
	.C(n_101), 
	.B(n_396), 
	.A(n_248));
   OA22X4 g28799 (.Q(n_544), 
	.D(n_186), 
	.C(n_98), 
	.B(n_394), 
	.A(n_154));
   AN22X2 g28800 (.Q(n_543), 
	.D(n_150), 
	.C(n_183), 
	.B(n_389), 
	.A(n_239));
   AN22X2 g28801 (.Q(n_542), 
	.D(n_119), 
	.C(n_279), 
	.B(n_406), 
	.A(n_90));
   AN21X4 g28802 (.Q(n_541), 
	.C(n_444), 
	.B(n_66), 
	.A(n_110));
   AN22X2 g28803 (.Q(n_540), 
	.D(n_288), 
	.C(n_96), 
	.B(n_390), 
	.A(n_68));
   OA22X4 g28804 (.Q(n_539), 
	.D(n_65), 
	.C(n_159), 
	.B(n_403), 
	.A(n_230));
   AN22X2 g28805 (.Q(n_538), 
	.D(n_126), 
	.C(n_3), 
	.B(n_393), 
	.A(n_269));
   AN22X2 g28806 (.Q(n_537), 
	.D(n_217), 
	.C(n_267), 
	.B(n_402), 
	.A(n_116));
   AN21X4 g28807 (.Q(n_536), 
	.C(n_446), 
	.B(n_88), 
	.A(n_40));
   AN21X4 g28808 (.Q(n_535), 
	.C(n_400), 
	.B(n_391), 
	.A(n_260));
   AN22X2 g28809 (.Q(n_534), 
	.D(n_123), 
	.C(n_66), 
	.B(n_404), 
	.A(n_321));
   OA22X4 g28810 (.Q(n_533), 
	.D(n_87), 
	.C(n_240), 
	.B(n_384), 
	.A(n_105));
   AN22X2 g28811 (.Q(n_532), 
	.D(n_71), 
	.C(n_183), 
	.B(n_389), 
	.A(n_283));
   AN22X2 g28812 (.Q(n_531), 
	.D(n_210), 
	.C(n_88), 
	.B(n_385), 
	.A(n_166));
   AN22X2 g28813 (.Q(n_530), 
	.D(n_222), 
	.C(n_183), 
	.B(n_389), 
	.A(n_281));
   OA22X4 g28814 (.Q(n_529), 
	.D(n_305), 
	.C(n_221), 
	.B(n_392), 
	.A(n_134));
   AN22X2 g28815 (.Q(n_528), 
	.D(n_119), 
	.C(n_62), 
	.B(n_406), 
	.A(n_273));
   AN22X2 g28816 (.Q(n_527), 
	.D(n_174), 
	.C(n_185), 
	.B(n_387), 
	.A(n_129));
   ON22X4 g28817 (.Q(n_526), 
	.D(n_118), 
	.C(n_103), 
	.B(n_405), 
	.A(n_202));
   AN22X2 g28818 (.Q(n_525), 
	.D(n_270), 
	.C(n_3), 
	.B(n_393), 
	.A(n_234));
   AO22X4 g28819 (.Q(n_524), 
	.D(n_183), 
	.C(n_281), 
	.B(n_389), 
	.A(n_115));
   AN21X2  g28820 (.Q(n_523), 
	.C(n_398), 
	.B(n_402), 
	.A(n_191));
   AN22X2 g28821 (.Q(n_522), 
	.D(n_183), 
	.C(n_239), 
	.B(n_389), 
	.A(n_70));
   AN22X2 g28822 (.Q(n_521), 
	.D(n_248), 
	.C(n_101), 
	.B(n_396), 
	.A(n_292));
   AN22X2 g28823 (.Q(n_520), 
	.D(n_116), 
	.C(n_267), 
	.B(n_402), 
	.A(n_249));
   AN22X2 g28824 (.Q(n_519), 
	.D(n_172), 
	.C(n_174), 
	.B(n_387), 
	.A(n_144));
   AN22X2 g28825 (.Q(n_518), 
	.D(n_292), 
	.C(n_101), 
	.B(n_396), 
	.A(n_137));
   AO22X4 g28826 (.Q(n_517), 
	.D(n_66), 
	.C(n_212), 
	.B(n_404), 
	.A(n_180));
   AN22X2 g28827 (.Q(n_516), 
	.D(n_227), 
	.C(n_101), 
	.B(n_396), 
	.A(n_86));
   ON22X4 g28828 (.Q(n_515), 
	.D(n_173), 
	.C(n_177), 
	.B(n_386), 
	.A(n_160));
   AN22X2 g28829 (.Q(n_514), 
	.D(n_267), 
	.C(n_249), 
	.B(n_402), 
	.A(n_42));
   AN22X2 g28830 (.Q(n_513), 
	.D(n_96), 
	.C(n_258), 
	.B(n_390), 
	.A(n_58));
   AN22X2 g28831 (.Q(n_512), 
	.D(n_231), 
	.C(n_3), 
	.B(n_393), 
	.A(n_57));
   OA22X4 g28832 (.Q(n_511), 
	.D(n_87), 
	.C(n_105), 
	.B(n_384), 
	.A(n_280));
   AN22X2 g28833 (.Q(n_510), 
	.D(n_68), 
	.C(n_96), 
	.B(n_390), 
	.A(n_245));
   AN22X2 g28834 (.Q(n_509), 
	.D(n_88), 
	.C(n_166), 
	.B(n_385), 
	.A(n_92));
   AO22X4 g28835 (.Q(n_508), 
	.D(n_119), 
	.C(n_257), 
	.B(n_406), 
	.A(n_287));
   AN22X2 g28836 (.Q(n_507), 
	.D(n_269), 
	.C(n_3), 
	.B(n_393), 
	.A(n_231));
   AN22X2 g28837 (.Q(n_506), 
	.D(n_272), 
	.C(n_304), 
	.B(n_391), 
	.A(n_247));
   AN22X2 g28838 (.Q(n_505), 
	.D(n_245), 
	.C(n_96), 
	.B(n_390), 
	.A(n_69));
   AO22X4 g28839 (.Q(n_504), 
	.D(n_267), 
	.C(n_218), 
	.B(n_402), 
	.A(n_78));
   AO22X4 g28840 (.Q(n_503), 
	.D(n_66), 
	.C(n_125), 
	.B(n_404), 
	.A(n_97));
   ON22X4 g28841 (.Q(n_502), 
	.D(n_186), 
	.C(n_47), 
	.B(n_394), 
	.A(n_82));
   OA22X4 g28842 (.Q(n_501), 
	.D(n_186), 
	.C(n_60), 
	.B(n_394), 
	.A(n_251));
   AN22X2 g28843 (.Q(n_500), 
	.D(n_225), 
	.C(n_101), 
	.B(n_396), 
	.A(n_161));
   AN22X2 g28844 (.Q(n_499), 
	.D(n_119), 
	.C(n_170), 
	.B(n_406), 
	.A(n_63));
   OA22X4 g28845 (.Q(n_498), 
	.D(n_100), 
	.C(n_142), 
	.B(n_395), 
	.A(n_213));
   AN22X2 g28846 (.Q(n_497), 
	.D(n_174), 
	.C(n_129), 
	.B(n_387), 
	.A(n_79));
   AN22X2 g28847 (.Q(n_496), 
	.D(n_83), 
	.C(n_66), 
	.B(n_404), 
	.A(n_49));
   ON22X4 g28848 (.Q(n_495), 
	.D(n_186), 
	.C(n_154), 
	.B(n_394), 
	.A(n_275));
   AN21X4 g28849 (.Q(n_494), 
	.C(n_445), 
	.B(n_3), 
	.A(n_57));
   AO22X4 g28850 (.Q(n_493), 
	.D(n_66), 
	.C(n_149), 
	.B(n_404), 
	.A(n_102));
   AN22X2 g28851 (.Q(n_492), 
	.D(n_267), 
	.C(n_42), 
	.B(n_402), 
	.A(n_53));
   AN22X2 g28852 (.Q(n_491), 
	.D(n_183), 
	.C(n_228), 
	.B(n_389), 
	.A(n_199));
   AN22X2 g28853 (.Q(n_490), 
	.D(n_164), 
	.C(n_96), 
	.B(n_390), 
	.A(n_89));
   AN22X2 g28854 (.Q(n_489), 
	.D(n_101), 
	.C(n_137), 
	.B(n_396), 
	.A(n_84));
   AN22X2 g28855 (.Q(n_488), 
	.D(n_101), 
	.C(n_84), 
	.B(n_396), 
	.A(n_233));
   ON22X4 g28856 (.Q(n_487), 
	.D(n_182), 
	.C(n_169), 
	.B(n_388), 
	.A(n_59));
   AN22X2 g28857 (.Q(n_486), 
	.D(n_183), 
	.C(n_199), 
	.B(n_389), 
	.A(n_318));
   AN22X2 g28858 (.Q(n_485), 
	.D(n_122), 
	.C(n_88), 
	.B(n_385), 
	.A(n_219));
   ON22X4 g28859 (.Q(n_484), 
	.D(n_100), 
	.C(n_213), 
	.B(n_395), 
	.A(n_139));
   AN22X2 g28860 (.Q(n_483), 
	.D(n_271), 
	.C(n_96), 
	.B(n_390), 
	.A(n_164));
   AN22X2 g28861 (.Q(n_482), 
	.D(n_250), 
	.C(n_96), 
	.B(n_390), 
	.A(n_51));
   AN22X2 g28862 (.Q(n_481), 
	.D(n_101), 
	.C(n_233), 
	.B(n_396), 
	.A(n_204));
   AN22X2 g28863 (.Q(n_480), 
	.D(n_119), 
	.C(n_287), 
	.B(n_406), 
	.A(n_133));
   OA22X4 g28864 (.Q(n_479), 
	.D(n_87), 
	.C(n_280), 
	.B(n_384), 
	.A(n_75));
   OA22X4 g28865 (.Q(n_478), 
	.D(n_186), 
	.C(n_179), 
	.B(n_394), 
	.A(n_95));
   AN21X4 g28866 (.Q(n_477), 
	.C(n_399), 
	.B(n_404), 
	.A(n_262));
   AN22X2 g28867 (.Q(n_476), 
	.D(n_267), 
	.C(n_226), 
	.B(n_402), 
	.A(n_327));
   ON22X4 g28868 (.Q(n_475), 
	.D(n_173), 
	.C(n_286), 
	.B(n_386), 
	.A(n_121));
   ON22X4 g28869 (.Q(n_474), 
	.D(n_186), 
	.C(n_82), 
	.B(n_394), 
	.A(n_45));
   AO22X4 g28870 (.Q(n_473), 
	.D(n_267), 
	.C(n_131), 
	.B(n_402), 
	.A(n_73));
   AN22X2 g28871 (.Q(n_472), 
	.D(n_72), 
	.C(n_304), 
	.B(n_391), 
	.A(n_254));
   AN22X2 g28872 (.Q(n_471), 
	.D(n_61), 
	.C(n_88), 
	.B(n_385), 
	.A(n_163));
   AN22X2 g28873 (.Q(n_470), 
	.D(n_101), 
	.C(n_204), 
	.B(n_396), 
	.A(n_54));
   AO22X4 g28874 (.Q(n_469), 
	.D(n_181), 
	.C(n_267), 
	.B(n_402), 
	.A(n_226));
   AN22X2 g28875 (.Q(n_468), 
	.D(n_268), 
	.C(n_101), 
	.B(n_396), 
	.A(n_227));
   AN22X2 g28876 (.Q(n_467), 
	.D(n_119), 
	.C(n_214), 
	.B(n_406), 
	.A(n_52));
   AN21X4 g28877 (.Q(n_466), 
	.C(n_443), 
	.B(n_304), 
	.A(n_254));
   AN22X2 g28878 (.Q(n_465), 
	.D(n_174), 
	.C(n_252), 
	.B(n_387), 
	.A(n_285));
   AN22X2 g28879 (.Q(n_464), 
	.D(n_54), 
	.C(n_101), 
	.B(n_396), 
	.A(n_268));
   AN22X2 g28880 (.Q(n_463), 
	.D(n_74), 
	.C(n_88), 
	.B(n_385), 
	.A(n_35));
   AN22X2 g28881 (.Q(n_462), 
	.D(n_238), 
	.C(n_174), 
	.B(n_387), 
	.A(n_278));
   AN22X2 g28882 (.Q(n_461), 
	.D(n_163), 
	.C(n_88), 
	.B(n_385), 
	.A(n_64));
   OA22X4 g28883 (.Q(n_460), 
	.D(n_186), 
	.C(n_95), 
	.B(n_394), 
	.A(n_232));
   AO22X4 g28884 (.Q(n_459), 
	.D(n_66), 
	.C(n_180), 
	.B(n_404), 
	.A(n_223));
   AN22X2 g28885 (.Q(n_458), 
	.D(n_229), 
	.C(n_66), 
	.B(n_404), 
	.A(n_125));
   NA2X4 g28886 (.Q(n_457), 
	.B(n_349), 
	.A(B[11]));
   NA2X4 g28887 (.Q(n_456), 
	.B(n_344), 
	.A(B[9]));
   NA2X4 g28888 (.Q(n_455), 
	.B(n_350), 
	.A(B[3]));
   NA2X4 g28889 (.Q(n_454), 
	.B(n_343), 
	.A(B[19]));
   NA2X4 g28890 (.Q(n_453), 
	.B(n_347), 
	.A(B[7]));
   NA2X4 g28891 (.Q(n_452), 
	.B(n_348), 
	.A(B[5]));
   NA2X4 g28892 (.Q(n_451), 
	.B(n_346), 
	.A(B[21]));
   NA2X4 g28893 (.Q(n_450), 
	.B(n_341), 
	.A(B[13]));
   NA2X4 g28894 (.Q(n_449), 
	.B(n_345), 
	.A(B[15]));
   NA2X4 g28895 (.Q(n_448), 
	.B(n_342), 
	.A(B[17]));
   NA2X4 g28896 (.Q(n_447), 
	.B(n_351), 
	.A(B[23]));
   NO2X4 g28897 (.Q(n_446), 
	.B(n_384), 
	.A(n_265));
   NO2X4 g28898 (.Q(n_445), 
	.B(n_394), 
	.A(n_60));
   NO2X4 g28899 (.Q(n_444), 
	.B(n_403), 
	.A(n_158));
   NO2X4 g28900 (.Q(n_443), 
	.B(n_392), 
	.A(n_221));
   AN22X2 g28901 (.Q(n_442), 
	.D(B[1]), 
	.C(B[0]), 
	.B(n_0), 
	.A(n_294));
   AN22X2 g28902 (.Q(n_441), 
	.D(n_303), 
	.C(B[0]), 
	.B(n_298), 
	.A(n_0));
   AN22X2 g28903 (.Q(n_440), 
	.D(B[0]), 
	.C(n_299), 
	.B(n_302), 
	.A(n_0));
   AN22X2 g28904 (.Q(n_439), 
	.D(n_307), 
	.C(B[0]), 
	.B(n_317), 
	.A(n_0));
   AN22X2 g28905 (.Q(n_438), 
	.D(B[0]), 
	.C(n_316), 
	.B(n_303), 
	.A(n_0));
   AN22X2 g28906 (.Q(n_437), 
	.D(n_302), 
	.C(B[0]), 
	.B(n_301), 
	.A(n_0));
   AN22X2 g28907 (.Q(n_436), 
	.D(n_301), 
	.C(B[0]), 
	.B(n_307), 
	.A(n_0));
   AN22X2 g28908 (.Q(n_435), 
	.D(n_313), 
	.C(B[0]), 
	.B(n_325), 
	.A(n_0));
   AN22X2 g28909 (.Q(n_434), 
	.D(n_309), 
	.C(B[0]), 
	.B(n_299), 
	.A(n_0));
   AN22X2 g28910 (.Q(n_433), 
	.D(n_310), 
	.C(B[0]), 
	.B(n_0), 
	.A(n_312));
   AN22X2 g28911 (.Q(n_432), 
	.D(n_298), 
	.C(B[0]), 
	.B(n_308), 
	.A(n_0));
   AN22X2 g28912 (.Q(n_431), 
	.D(n_312), 
	.C(B[0]), 
	.B(n_0), 
	.A(n_295));
   AN22X2 g28913 (.Q(n_430), 
	.D(n_306), 
	.C(B[0]), 
	.B(n_300), 
	.A(n_0));
   AN22X2 g28914 (.Q(n_429), 
	.D(B[0]), 
	.C(n_295), 
	.B(n_306), 
	.A(n_0));
   AN22X2 g28915 (.Q(n_428), 
	.D(n_297), 
	.C(B[0]), 
	.B(n_315), 
	.A(n_0));
   AN22X2 g28916 (.Q(n_427), 
	.D(B[0]), 
	.C(n_300), 
	.B(n_311), 
	.A(n_0));
   AN22X2 g28917 (.Q(n_426), 
	.D(B[0]), 
	.C(n_296), 
	.B(n_297), 
	.A(n_0));
   AN22X2 g28918 (.Q(n_425), 
	.D(n_311), 
	.C(B[0]), 
	.B(n_296), 
	.A(n_0));
   AN22X2 g28919 (.Q(n_424), 
	.D(B[0]), 
	.C(n_294), 
	.B(n_0), 
	.A(n_310));
   AN22X2 g28920 (.Q(n_423), 
	.D(B[0]), 
	.C(n_317), 
	.B(n_313), 
	.A(n_0));
   AN22X2 g28921 (.Q(n_422), 
	.D(n_308), 
	.C(B[0]), 
	.B(n_309), 
	.A(n_0));
   AN22X2 g28922 (.Q(n_421), 
	.D(B[0]), 
	.C(n_315), 
	.B(n_293), 
	.A(n_0));
   AN22X2 g28923 (.Q(n_420), 
	.D(n_293), 
	.C(B[0]), 
	.B(n_314), 
	.A(n_0));
   AN22X2 g28924 (.Q(n_419), 
	.D(B[0]), 
	.C(n_314), 
	.B(n_316), 
	.A(n_0));
   NA2X4 g28925 (.Q(n_418), 
	.B(n_183), 
	.A(A[0]));
   NA2X4 g28926 (.Q(n_417), 
	.B(n_304), 
	.A(A[0]));
   NA2X4 g28927 (.Q(n_416), 
	.B(n_174), 
	.A(A[0]));
   NA2X4 g28928 (.Q(n_415), 
	.B(n_2), 
	.A(A[0]));
   NA2X4 g28929 (.Q(n_414), 
	.B(n_66), 
	.A(A[0]));
   NA2X4 g28930 (.Q(n_413), 
	.B(n_119), 
	.A(A[0]));
   NA2X4 g28931 (.Q(n_412), 
	.B(n_267), 
	.A(A[0]));
   NA2X4 g28932 (.Q(n_411), 
	.B(n_3), 
	.A(A[0]));
   NA2X4 g28933 (.Q(n_410), 
	.B(n_101), 
	.A(A[0]));
   NA2X4 g28934 (.Q(n_409), 
	.B(n_88), 
	.A(A[0]));
   NA2X4 g28935 (.Q(n_408), 
	.B(n_96), 
	.A(A[0]));
   NO2X4 g28936 (.Q(n_407), 
	.B(n_305), 
	.A(n_187));
   INX8 g28937 (.Q(n_405), 
	.A(n_406));
   NO2X4 g28938 (.Q(n_406), 
	.B(n_119), 
	.A(n_335));
   INX8 g28939 (.Q(n_403), 
	.A(n_404));
   NO2X3 g28940 (.Q(n_404), 
	.B(n_66), 
	.A(n_339));
   INX8 g28941 (.Q(n_401), 
	.A(n_402));
   NO2X4 g28942 (.Q(n_402), 
	.B(n_267), 
	.A(n_336));
   NO2X4 g28943 (.Q(n_400), 
	.B(n_305), 
	.A(n_108));
   NO2X4 g28944 (.Q(n_399), 
	.B(n_65), 
	.A(n_143));
   NO2X4 g28945 (.Q(n_398), 
	.B(n_266), 
	.A(n_148));
   NO2X4 g28946 (.Q(n_397), 
	.B(n_2), 
	.A(n_334));
   INX8 g28947 (.Q(n_395), 
	.A(n_396));
   AND2X4 g28948 (.Q(n_396), 
	.B(n_100), 
	.A(n_337));
   INX8 g28949 (.Q(n_393), 
	.A(n_394));
   OR2X3 g28950 (.Q(n_394), 
	.B(n_3), 
	.A(n_329));
   INX8 g28951 (.Q(n_391), 
	.A(n_392));
   OR2X4 g28952 (.Q(n_392), 
	.B(n_304), 
	.A(n_332));
   NO2X4 g28953 (.Q(n_390), 
	.B(n_96), 
	.A(n_330));
   INX8 g28954 (.Q(n_388), 
	.A(n_389));
   AND2X4 g28955 (.Q(n_389), 
	.B(n_182), 
	.A(n_338));
   INX8 g28956 (.Q(n_386), 
	.A(n_387));
   NO2X3 g28957 (.Q(n_387), 
	.B(n_174), 
	.A(n_331));
   INX8 g28958 (.Q(n_384), 
	.A(n_385));
   AND2X4 g28959 (.Q(n_385), 
	.B(n_87), 
	.A(n_333));
   HAX4 g28960 (.S(n_383), 
	.CO(n_382), 
	.B(A[11]), 
	.A(B[23]));
   HAX4 g28961 (.S(n_380), 
	.CO(n_381), 
	.B(A[0]), 
	.A(B[23]));
   HAX4 g28962 (.S(n_379), 
	.CO(n_378), 
	.B(A[19]), 
	.A(B[23]));
   HAX4 g28963 (.S(n_377), 
	.CO(n_376), 
	.B(A[6]), 
	.A(B[23]));
   HAX4 g28964 (.S(n_375), 
	.CO(n_374), 
	.B(A[3]), 
	.A(B[23]));
   HAX4 g28965 (.S(n_373), 
	.CO(n_372), 
	.B(A[20]), 
	.A(B[23]));
   HAX4 g28966 (.S(n_371), 
	.CO(n_370), 
	.B(A[18]), 
	.A(B[23]));
   HAX4 g28967 (.S(n_369), 
	.CO(n_368), 
	.B(A[7]), 
	.A(B[23]));
   HAX4 g28968 (.S(n_367), 
	.CO(n_366), 
	.B(A[17]), 
	.A(B[23]));
   HAX4 g28969 (.S(n_365), 
	.CO(n_364), 
	.B(A[21]), 
	.A(B[23]));
   HAX4 g28970 (.S(n_363), 
	.CO(n_362), 
	.B(A[8]), 
	.A(B[23]));
   HAX4 g28971 (.S(n_361), 
	.CO(n_360), 
	.B(A[23]), 
	.A(B[23]));
   HAX4 g28972 (.S(n_359), 
	.CO(n_358), 
	.B(A[5]), 
	.A(B[23]));
   HAX4 g28973 (.S(n_357), 
	.CO(n_356), 
	.B(A[14]), 
	.A(B[23]));
   HAX4 g28974 (.S(n_355), 
	.CO(n_354), 
	.B(A[2]), 
	.A(B[23]));
   HAX4 g28975 (.S(n_353), 
	.CO(n_352), 
	.B(A[22]), 
	.A(B[23]));
   EN3X2 g28976 (.Q(n_351), 
	.C(B[21]), 
	.B(B[22]), 
	.A(A[0]));
   EN3X2 g28977 (.Q(n_350), 
	.C(B[1]), 
	.B(B[2]), 
	.A(A[0]));
   EN3X2 g28978 (.Q(n_349), 
	.C(B[9]), 
	.B(B[10]), 
	.A(A[0]));
   EN3X2 g28979 (.Q(n_348), 
	.C(B[3]), 
	.B(B[4]), 
	.A(A[0]));
   EN3X2 g28980 (.Q(n_347), 
	.C(B[5]), 
	.B(B[6]), 
	.A(A[0]));
   EN3X2 g28981 (.Q(n_346), 
	.C(B[19]), 
	.B(B[20]), 
	.A(A[0]));
   EN3X2 g28982 (.Q(n_345), 
	.C(B[13]), 
	.B(B[14]), 
	.A(A[0]));
   EN3X2 g28983 (.Q(n_344), 
	.C(B[7]), 
	.B(B[8]), 
	.A(A[0]));
   EN3X2 g28984 (.Q(n_343), 
	.C(B[17]), 
	.B(B[18]), 
	.A(A[0]));
   EN3X2 g28985 (.Q(n_342), 
	.C(B[15]), 
	.B(B[16]), 
	.A(A[0]));
   EN3X2 g28986 (.Q(n_341), 
	.C(B[11]), 
	.B(B[12]), 
	.A(A[0]));
   NA2I1X4 g28987 (.Q(n_340), 
	.B(B[1]), 
	.AN(Z[0]));
   EN2X4 g28988 (.Q(n_339), 
	.B(B[19]), 
	.A(B[18]));
   EO2X3 g28989 (.Q(n_338), 
	.B(B[15]), 
	.A(B[14]));
   EO2X3 g28990 (.Q(n_337), 
	.B(B[7]), 
	.A(B[6]));
   EN2X4 g28991 (.Q(n_336), 
	.B(B[13]), 
	.A(B[12]));
   EN2X4 g28992 (.Q(n_335), 
	.B(B[17]), 
	.A(B[16]));
   EN2X4 g28993 (.Q(n_334), 
	.B(B[23]), 
	.A(B[22]));
   EO2X3 g28994 (.Q(n_333), 
	.B(B[9]), 
	.A(B[8]));
   EN2X4 g28995 (.Q(n_332), 
	.B(B[3]), 
	.A(B[2]));
   EN2X4 g28996 (.Q(n_331), 
	.B(B[21]), 
	.A(B[20]));
   EN2X4 g28997 (.Q(n_330), 
	.B(B[5]), 
	.A(B[4]));
   EN2X4 g28998 (.Q(n_329), 
	.B(B[11]), 
	.A(B[10]));
   EO2X3 g28999 (.Q(n_328), 
	.B(B[9]), 
	.A(A[0]));
   EO2X3 g29000 (.Q(n_327), 
	.B(B[13]), 
	.A(A[0]));
   EO2X3 g29001 (.Q(n_326), 
	.B(B[3]), 
	.A(A[0]));
   EO2X3 g29002 (.Q(n_325), 
	.B(B[1]), 
	.A(A[0]));
   EO2X3 g29003 (.Q(n_324), 
	.B(B[5]), 
	.A(A[0]));
   EO2X3 g29004 (.Q(n_323), 
	.B(B[21]), 
	.A(A[0]));
   EN2X4 g29005 (.Q(n_322), 
	.B(B[11]), 
	.A(A[0]));
   EO2X3 g29006 (.Q(n_321), 
	.B(B[19]), 
	.A(A[0]));
   EN2X4 g29007 (.Q(n_320), 
	.B(n_15), 
	.A(A[0]));
   EO2X3 g29008 (.Q(n_319), 
	.B(B[17]), 
	.A(A[0]));
   EO2X3 g29009 (.Q(n_318), 
	.B(B[15]), 
	.A(A[0]));
   EO2X3 g29010 (.Q(n_317), 
	.B(B[1]), 
	.A(A[2]));
   EO2X3 g29011 (.Q(n_316), 
	.B(B[1]), 
	.A(A[11]));
   EO2X3 g29012 (.Q(n_315), 
	.B(B[1]), 
	.A(A[14]));
   EO2X3 g29013 (.Q(n_314), 
	.B(B[1]), 
	.A(A[12]));
   EO2X3 g29014 (.Q(n_313), 
	.B(B[1]), 
	.A(A[1]));
   EO2X3 g29015 (.Q(n_312), 
	.B(B[1]), 
	.A(A[21]));
   EO2X3 g29016 (.Q(n_311), 
	.B(B[1]), 
	.A(A[17]));
   EO2X3 g29017 (.Q(n_310), 
	.B(B[1]), 
	.A(A[22]));
   EO2X3 g29018 (.Q(n_309), 
	.B(B[1]), 
	.A(A[7]));
   EO2X3 g29019 (.Q(n_308), 
	.B(B[1]), 
	.A(A[8]));
   EO2X3 g29020 (.Q(n_307), 
	.B(B[1]), 
	.A(A[3]));
   EO2X3 g29021 (.Q(n_306), 
	.B(B[1]), 
	.A(A[19]));
   INX8 g29022 (.Q(n_304), 
	.A(n_305));
   EN2X4 g29023 (.Q(n_305), 
	.B(B[1]), 
	.A(B[2]));
   EO2X3 g29024 (.Q(n_303), 
	.B(B[1]), 
	.A(A[10]));
   EO2X3 g29025 (.Q(n_302), 
	.B(B[1]), 
	.A(A[5]));
   EO2X3 g29026 (.Q(n_301), 
	.B(B[1]), 
	.A(A[4]));
   EO2X3 g29027 (.Q(n_300), 
	.B(B[1]), 
	.A(A[18]));
   EO2X3 g29028 (.Q(n_299), 
	.B(B[1]), 
	.A(A[6]));
   EO2X3 g29029 (.Q(n_298), 
	.B(B[1]), 
	.A(A[9]));
   EO2X3 g29030 (.Q(n_297), 
	.B(B[1]), 
	.A(A[15]));
   EO2X3 g29031 (.Q(n_296), 
	.B(B[1]), 
	.A(A[16]));
   EO2X3 g29032 (.Q(n_295), 
	.B(B[1]), 
	.A(A[20]));
   EO2X3 g29033 (.Q(n_294), 
	.B(B[1]), 
	.A(A[23]));
   EO2X3 g29034 (.Q(n_293), 
	.B(B[1]), 
	.A(A[13]));
   EO2X3 g29035 (.Q(n_292), 
	.B(B[7]), 
	.A(A[11]));
   EN2X4 g29036 (.Q(n_291), 
	.B(B[7]), 
	.A(A[23]));
   EO2X3 g29037 (.Q(n_290), 
	.B(B[13]), 
	.A(A[18]));
   EN2X4 g29038 (.Q(n_289), 
	.B(B[3]), 
	.A(A[22]));
   EO2X3 g29039 (.Q(n_288), 
	.B(B[5]), 
	.A(A[15]));
   EO2X3 g29040 (.Q(n_287), 
	.B(B[17]), 
	.A(A[10]));
   EN2X4 g29041 (.Q(n_286), 
	.B(B[21]), 
	.A(A[21]));
   EO2X3 g29042 (.Q(n_285), 
	.B(B[21]), 
	.A(A[4]));
   EO2X3 g29043 (.Q(n_284), 
	.B(B[9]), 
	.A(A[12]));
   INX4 g29044 (.Q(n_283), 
	.A(n_282));
   EN2X4 g29045 (.Q(n_282), 
	.B(B[15]), 
	.A(A[19]));
   EO2X3 g29046 (.Q(n_281), 
	.B(B[15]), 
	.A(A[13]));
   EN2X4 g29047 (.Q(n_280), 
	.B(B[9]), 
	.A(A[18]));
   EO2X3 g29048 (.Q(n_279), 
	.B(B[17]), 
	.A(A[8]));
   INX4 g29049 (.Q(n_278), 
	.A(n_277));
   EN2X4 g29050 (.Q(n_277), 
	.B(B[21]), 
	.A(A[12]));
   EO2X3 g29051 (.Q(n_276), 
	.B(B[5]), 
	.A(A[21]));
   INX4 g29052 (.Q(n_275), 
	.A(n_274));
   EO2X3 g29053 (.Q(n_274), 
	.B(B[11]), 
	.A(A[16]));
   EO2X3 g29054 (.Q(n_273), 
	.B(B[17]), 
	.A(A[21]));
   EO2X3 g29055 (.Q(n_272), 
	.B(B[3]), 
	.A(A[15]));
   EO2X3 g29056 (.Q(n_271), 
	.B(B[5]), 
	.A(A[19]));
   EO2X3 g29057 (.Q(n_270), 
	.B(B[11]), 
	.A(A[14]));
   EO2X3 g29058 (.Q(n_269), 
	.B(B[11]), 
	.A(A[8]));
   EO2X3 g29059 (.Q(n_268), 
	.B(B[7]), 
	.A(A[5]));
   INX8 g29060 (.Q(n_266), 
	.A(n_267));
   EN2X4 g29061 (.Q(n_267), 
	.B(n_17), 
	.A(B[12]));
   EN2X4 g29062 (.Q(n_265), 
	.B(B[9]), 
	.A(A[22]));
   EO2X3 g29063 (.Q(n_264), 
	.B(B[19]), 
	.A(A[4]));
   EN2X4 g29064 (.Q(n_263), 
	.B(B[3]), 
	.A(A[6]));
   EO2X3 g29065 (.Q(n_262), 
	.B(B[19]), 
	.A(A[7]));
   EO2X3 g29066 (.Q(n_261), 
	.B(B[9]), 
	.A(A[15]));
   EO2X3 g29067 (.Q(n_260), 
	.B(B[3]), 
	.A(A[16]));
   EO2X3 g29068 (.Q(n_259), 
	.B(B[11]), 
	.A(A[15]));
   EO2X3 g29069 (.Q(n_258), 
	.B(B[5]), 
	.A(A[23]));
   EO2X3 g29070 (.Q(n_257), 
	.B(B[17]), 
	.A(A[11]));
   EO2X3 g29071 (.Q(n_256), 
	.B(B[7]), 
	.A(A[18]));
   EO2X3 g29072 (.Q(n_255), 
	.B(B[7]), 
	.A(A[1]));
   EO2X3 g29073 (.Q(n_254), 
	.B(B[3]), 
	.A(A[10]));
   EO2X3 g29074 (.Q(n_253), 
	.B(B[5]), 
	.A(A[1]));
   EO2X3 g29075 (.Q(n_252), 
	.B(B[21]), 
	.A(A[5]));
   EN2X4 g29076 (.Q(n_251), 
	.B(B[11]), 
	.A(A[4]));
   EO2X3 g29077 (.Q(n_250), 
	.B(B[5]), 
	.A(A[10]));
   EO2X3 g29078 (.Q(n_249), 
	.B(B[13]), 
	.A(A[5]));
   EO2X3 g29079 (.Q(n_248), 
	.B(B[7]), 
	.A(A[12]));
   EO2X3 g29080 (.Q(n_247), 
	.B(B[3]), 
	.A(A[14]));
   EO2X3 g29081 (.Q(n_246), 
	.B(B[17]), 
	.A(A[23]));
   EO2X3 g29082 (.Q(n_245), 
	.B(B[5]), 
	.A(A[13]));
   EO2X3 g29083 (.Q(n_244), 
	.B(B[5]), 
	.A(A[3]));
   EO2X3 g29084 (.Q(n_243), 
	.B(B[17]), 
	.A(A[20]));
   EO2X3 g29085 (.Q(n_242), 
	.B(B[17]), 
	.A(A[19]));
   EO2X3 g29086 (.Q(n_241), 
	.B(B[17]), 
	.A(A[4]));
   EN2X4 g29087 (.Q(n_240), 
	.B(B[9]), 
	.A(A[20]));
   EO2X3 g29088 (.Q(n_239), 
	.B(B[15]), 
	.A(A[4]));
   EO2X3 g29089 (.Q(n_238), 
	.B(B[21]), 
	.A(A[13]));
   EO2X3 g29090 (.Q(n_237), 
	.B(B[21]), 
	.A(A[3]));
   EO2X3 g29091 (.Q(n_236), 
	.B(B[21]), 
	.A(A[9]));
   EO2X3 g29092 (.Q(n_235), 
	.B(B[3]), 
	.A(A[12]));
   EO2X3 g29093 (.Q(n_234), 
	.B(B[11]), 
	.A(A[13]));
   EO2X3 g29094 (.Q(n_233), 
	.B(B[7]), 
	.A(A[8]));
   EN2X4 g29095 (.Q(n_232), 
	.B(B[11]), 
	.A(A[1]));
   EO2X3 g29096 (.Q(n_231), 
	.B(B[11]), 
	.A(A[7]));
   INX4 g29097 (.Q(n_230), 
	.A(n_229));
   EO2X3 g29098 (.Q(n_229), 
	.B(B[19]), 
	.A(A[15]));
   EO2X3 g29099 (.Q(n_228), 
	.B(B[15]), 
	.A(A[2]));
   EO2X3 g29100 (.Q(n_227), 
	.B(B[7]), 
	.A(A[4]));
   EO2X3 g29101 (.Q(n_226), 
	.B(B[13]), 
	.A(A[1]));
   EO2X3 g29102 (.Q(n_225), 
	.B(B[7]), 
	.A(A[17]));
   EO2X3 g29103 (.Q(n_224), 
	.B(B[5]), 
	.A(A[5]));
   EO2X3 g29104 (.Q(n_223), 
	.B(B[19]), 
	.A(A[21]));
   EO2X3 g29105 (.Q(n_222), 
	.B(B[15]), 
	.A(A[14]));
   EN2X4 g29106 (.Q(n_221), 
	.B(B[3]), 
	.A(A[9]));
   EO2X3 g29107 (.Q(n_220), 
	.B(B[17]), 
	.A(A[3]));
   EO2X3 g29108 (.Q(n_219), 
	.B(B[9]), 
	.A(A[6]));
   EO2X3 g29109 (.Q(n_218), 
	.B(B[13]), 
	.A(A[15]));
   EO2X3 g29110 (.Q(n_217), 
	.B(B[13]), 
	.A(A[7]));
   EO2X3 g29111 (.Q(n_216), 
	.B(B[5]), 
	.A(A[16]));
   EO2X3 g29112 (.Q(n_215), 
	.B(B[13]), 
	.A(A[11]));
   EO2X3 g29113 (.Q(n_214), 
	.B(B[17]), 
	.A(A[6]));
   EN2X4 g29114 (.Q(n_213), 
	.B(B[7]), 
	.A(A[20]));
   EO2X3 g29115 (.Q(n_212), 
	.B(B[19]), 
	.A(A[23]));
   EO2X3 g29116 (.Q(n_211), 
	.B(B[15]), 
	.A(A[9]));
   EO2X3 g29117 (.Q(n_210), 
	.B(B[9]), 
	.A(A[11]));
   EN2X4 g29118 (.Q(n_209), 
	.B(B[3]), 
	.A(A[20]));
   EO2X3 g29119 (.Q(n_208), 
	.B(B[13]), 
	.A(A[17]));
   EN2X4 g29120 (.Q(n_207), 
	.B(B[3]), 
	.A(A[21]));
   EO2X3 g29121 (.Q(n_206), 
	.B(B[5]), 
	.A(A[2]));
   EO2X3 g29122 (.Q(n_205), 
	.B(B[15]), 
	.A(A[8]));
   EO2X3 g29123 (.Q(n_204), 
	.B(B[7]), 
	.A(A[7]));
   EO2X3 g29124 (.Q(n_203), 
	.B(B[21]), 
	.A(A[2]));
   EN2X4 g29125 (.Q(n_202), 
	.B(B[17]), 
	.A(A[15]));
   EO2X3 g29126 (.Q(n_201), 
	.B(B[19]), 
	.A(A[12]));
   EO2X3 g29127 (.Q(n_200), 
	.B(B[9]), 
	.A(A[14]));
   EO2X3 g29128 (.Q(n_199), 
	.B(B[15]), 
	.A(A[1]));
   EO2X3 g29129 (.Q(n_198), 
	.B(B[7]), 
	.A(A[13]));
   EO2X3 g29130 (.Q(n_197), 
	.B(B[11]), 
	.A(A[12]));
   EN2X4 g29131 (.Q(n_196), 
	.B(B[11]), 
	.A(A[19]));
   EN2X4 g29132 (.Q(n_195), 
	.B(B[3]), 
	.A(A[4]));
   EN2X4 g29133 (.Q(n_194), 
	.B(B[3]), 
	.A(A[19]));
   EO2X3 g29134 (.Q(n_193), 
	.B(B[19]), 
	.A(A[3]));
   EN2X4 g29135 (.Q(n_192), 
	.B(B[9]), 
	.A(A[21]));
   EO2X3 g29136 (.Q(n_191), 
	.B(B[13]), 
	.A(A[21]));
   EO2X3 g29137 (.Q(n_190), 
	.B(B[11]), 
	.A(A[11]));
   EO2X3 g29138 (.Q(n_189), 
	.B(B[15]), 
	.A(A[21]));
   EN2X4 g29139 (.Q(n_188), 
	.B(B[3]), 
	.A(A[18]));
   EN2X4 g29140 (.Q(n_187), 
	.B(B[3]), 
	.A(A[3]));
   INX8 g29141 (.Q(n_186), 
	.A(n_3));
   EO2X3 g29143 (.Q(n_185), 
	.B(B[21]), 
	.A(A[8]));
   EO2X3 g29144 (.Q(n_184), 
	.B(B[21]), 
	.A(A[15]));
   INX8 g29145 (.Q(n_182), 
	.A(n_183));
   EN2X4 g29146 (.Q(n_183), 
	.B(n_13), 
	.A(B[14]));
   EO2X3 g29147 (.Q(n_181), 
	.B(B[13]), 
	.A(A[2]));
   EO2X3 g29148 (.Q(n_180), 
	.B(B[19]), 
	.A(A[22]));
   EN2X4 g29149 (.Q(n_179), 
	.B(B[11]), 
	.A(A[3]));
   INX4 g29150 (.Q(n_178), 
	.A(n_177));
   EN2X4 g29151 (.Q(n_177), 
	.B(B[21]), 
	.A(A[23]));
   EO2X3 g29152 (.Q(n_176), 
	.B(B[5]), 
	.A(A[4]));
   EO2X3 g29153 (.Q(n_175), 
	.B(B[15]), 
	.A(A[7]));
   INX8 g29154 (.Q(n_173), 
	.A(n_174));
   EO2X3 g29155 (.Q(n_174), 
	.B(B[20]), 
	.A(B[19]));
   EO2X3 g29156 (.Q(n_172), 
	.B(B[21]), 
	.A(A[19]));
   EO2X3 g29157 (.Q(n_171), 
	.B(B[5]), 
	.A(A[20]));
   EO2X3 g29158 (.Q(n_170), 
	.B(B[17]), 
	.A(A[18]));
   EN2X4 g29159 (.Q(n_169), 
	.B(B[15]), 
	.A(A[18]));
   EO2X3 g29160 (.Q(n_168), 
	.B(B[11]), 
	.A(A[10]));
   EO2X3 g29161 (.Q(n_167), 
	.B(B[5]), 
	.A(A[8]));
   EO2X3 g29162 (.Q(n_166), 
	.B(B[9]), 
	.A(A[10]));
   EO2X3 g29163 (.Q(n_165), 
	.B(B[13]), 
	.A(A[9]));
   EO2X3 g29164 (.Q(n_164), 
	.B(B[5]), 
	.A(A[18]));
   EO2X3 g29165 (.Q(n_163), 
	.B(B[9]), 
	.A(A[4]));
   EN2X4 g29166 (.Q(n_162), 
	.B(n_14), 
	.A(A[1]));
   EO2X3 g29167 (.Q(n_161), 
	.B(B[7]), 
	.A(A[16]));
   EN2X4 g29168 (.Q(n_160), 
	.B(B[21]), 
	.A(A[22]));
   EN2X4 g29169 (.Q(n_159), 
	.B(B[19]), 
	.A(A[16]));
   EN2X4 g29170 (.Q(n_158), 
	.B(B[19]), 
	.A(A[9]));
   EO2X3 g29171 (.Q(n_157), 
	.B(B[15]), 
	.A(A[6]));
   EO2X3 g29172 (.Q(n_156), 
	.B(B[13]), 
	.A(A[8]));
   EO2X3 g29173 (.Q(n_155), 
	.B(B[3]), 
	.A(A[13]));
   EN2X4 g29174 (.Q(n_154), 
	.B(B[11]), 
	.A(A[17]));
   EO2X3 g29175 (.Q(n_153), 
	.B(B[21]), 
	.A(A[17]));
   EO2X3 g29176 (.Q(n_152), 
	.B(B[13]), 
	.A(A[12]));
   EO2X3 g29177 (.Q(n_151), 
	.B(B[5]), 
	.A(A[6]));
   EO2X3 g29178 (.Q(n_150), 
	.B(B[15]), 
	.A(A[5]));
   EO2X3 g29179 (.Q(n_149), 
	.B(B[19]), 
	.A(A[20]));
   EN2X4 g29180 (.Q(n_148), 
	.B(B[13]), 
	.A(A[22]));
   EO2X3 g29181 (.Q(n_147), 
	.B(B[13]), 
	.A(A[13]));
   EO2X3 g29182 (.Q(n_146), 
	.B(B[3]), 
	.A(A[2]));
   EO2X3 g29183 (.Q(n_145), 
	.B(B[15]), 
	.A(A[22]));
   EO2X3 g29184 (.Q(n_144), 
	.B(B[21]), 
	.A(A[18]));
   EN2X4 g29185 (.Q(n_143), 
	.B(B[19]), 
	.A(A[8]));
   EN2X4 g29186 (.Q(n_142), 
	.B(B[7]), 
	.A(A[21]));
   EO2X3 g29187 (.Q(n_141), 
	.B(B[21]), 
	.A(A[16]));
   EO2X3 g29188 (.Q(n_140), 
	.B(B[17]), 
	.A(A[12]));
   INX4 g29189 (.Q(n_139), 
	.A(n_138));
   EO2X3 g29190 (.Q(n_138), 
	.B(B[7]), 
	.A(A[19]));
   EO2X3 g29191 (.Q(n_137), 
	.B(B[7]), 
	.A(A[10]));
   EN2X4 g29192 (.Q(n_136), 
	.B(B[17]), 
	.A(A[14]));
   EO2X3 g29193 (.Q(n_135), 
	.B(B[7]), 
	.A(A[15]));
   EN2X4 g29194 (.Q(n_134), 
	.B(B[3]), 
	.A(A[8]));
   EO2X3 g29195 (.Q(n_133), 
	.B(B[17]), 
	.A(A[9]));
   EO2X3 g29196 (.Q(n_132), 
	.B(B[19]), 
	.A(A[6]));
   EO2X3 g29197 (.Q(n_131), 
	.B(B[13]), 
	.A(A[20]));
   EO2X3 g29198 (.Q(n_130), 
	.B(B[17]), 
	.A(A[2]));
   EO2X3 g29199 (.Q(n_129), 
	.B(B[21]), 
	.A(A[7]));
   EO2X3 g29200 (.Q(n_128), 
	.B(B[15]), 
	.A(A[10]));
   EO2X3 g29201 (.Q(n_127), 
	.B(B[21]), 
	.A(A[1]));
   EO2X3 g29202 (.Q(n_126), 
	.B(B[11]), 
	.A(A[9]));
   EO2X3 g29203 (.Q(n_125), 
	.B(B[19]), 
	.A(A[14]));
   EN2X4 g29204 (.Q(n_124), 
	.B(B[15]), 
	.A(A[16]));
   EO2X3 g29205 (.Q(n_123), 
	.B(B[19]), 
	.A(A[1]));
   EO2X3 g29206 (.Q(n_122), 
	.B(B[9]), 
	.A(A[7]));
   INX4 g29207 (.Q(n_121), 
	.A(n_120));
   EO2X3 g29208 (.Q(n_120), 
	.B(B[21]), 
	.A(A[20]));
   INX8 g29209 (.Q(n_118), 
	.A(n_119));
   EN2X4 g29210 (.Q(n_119), 
	.B(n_16), 
	.A(B[16]));
   EO2X3 g29211 (.Q(n_117), 
	.B(B[19]), 
	.A(A[5]));
   EO2X3 g29212 (.Q(n_116), 
	.B(B[13]), 
	.A(A[6]));
   EO2X3 g29213 (.Q(n_115), 
	.B(B[15]), 
	.A(A[12]));
   EN2X4 g29214 (.Q(n_114), 
	.B(B[11]), 
	.A(A[20]));
   EO2X3 g29215 (.Q(n_113), 
	.B(B[19]), 
	.A(A[2]));
   INX4 g29216 (.Q(n_112), 
	.A(n_111));
   EO2X3 g29217 (.Q(n_111), 
	.B(B[21]), 
	.A(A[10]));
   EO2X3 g29218 (.Q(n_110), 
	.B(B[19]), 
	.A(A[10]));
   EO2X3 g29219 (.Q(n_109), 
	.B(B[17]), 
	.A(A[1]));
   EN2X4 g29220 (.Q(n_108), 
	.B(B[3]), 
	.A(A[17]));
   EO2X3 g29221 (.Q(n_107), 
	.B(B[19]), 
	.A(A[11]));
   EN2X4 g29222 (.Q(n_106), 
	.B(B[3]), 
	.A(A[23]));
   EN2X4 g29223 (.Q(n_105), 
	.B(B[9]), 
	.A(A[19]));
   INX4 g29224 (.Q(n_104), 
	.A(n_103));
   EN2X4 g29225 (.Q(n_103), 
	.B(B[17]), 
	.A(A[16]));
   EO2X3 g29226 (.Q(n_102), 
	.B(B[19]), 
	.A(A[19]));
   INX8 g29227 (.Q(n_100), 
	.A(n_101));
   EO2X3 g29228 (.Q(n_101), 
	.B(B[6]), 
	.A(B[5]));
   EO2X3 g29229 (.Q(n_99), 
	.B(B[5]), 
	.A(A[7]));
   EN2X4 g29230 (.Q(n_98), 
	.B(B[11]), 
	.A(A[18]));
   EO2X3 g29231 (.Q(n_97), 
	.B(B[19]), 
	.A(A[13]));
   EN2X4 g29232 (.Q(n_96), 
	.B(n_14), 
	.A(B[4]));
   EN2X4 g29233 (.Q(n_95), 
	.B(B[11]), 
	.A(A[2]));
   EO2X3 g29234 (.Q(n_94), 
	.B(B[21]), 
	.A(A[14]));
   EO2X3 g29235 (.Q(n_93), 
	.B(B[7]), 
	.A(A[2]));
   EO2X3 g29236 (.Q(n_92), 
	.B(B[9]), 
	.A(A[9]));
   EO2X3 g29237 (.Q(n_91), 
	.B(B[9]), 
	.A(A[13]));
   EO2X3 g29238 (.Q(n_90), 
	.B(B[17]), 
	.A(A[7]));
   EO2X3 g29239 (.Q(n_89), 
	.B(B[5]), 
	.A(A[17]));
   INX8 g29240 (.Q(n_87), 
	.A(n_88));
   EN2X4 g29241 (.Q(n_88), 
	.B(n_15), 
	.A(B[8]));
   EO2X3 g29242 (.Q(n_86), 
	.B(B[7]), 
	.A(A[3]));
   EO2X3 g29243 (.Q(n_85), 
	.B(B[9]), 
	.A(A[8]));
   EO2X3 g29244 (.Q(n_84), 
	.B(B[7]), 
	.A(A[9]));
   EO2X3 g29245 (.Q(n_83), 
	.B(B[19]), 
	.A(A[18]));
   EN2X4 g29246 (.Q(n_82), 
	.B(B[11]), 
	.A(A[22]));
   EO2X3 g29247 (.Q(n_81), 
	.B(B[9]), 
	.A(A[2]));
   EO2X3 g29248 (.Q(n_80), 
	.B(B[5]), 
	.A(A[11]));
   EO2X3 g29249 (.Q(n_79), 
	.B(B[21]), 
	.A(A[6]));
   EO2X3 g29250 (.Q(n_78), 
	.B(B[13]), 
	.A(A[14]));
   EO2X3 g29251 (.Q(n_77), 
	.B(B[15]), 
	.A(A[23]));
   EN2X4 g29252 (.Q(n_76), 
	.B(B[13]), 
	.A(A[23]));
   INX4 g29253 (.Q(n_75), 
	.A(n_74));
   EO2X3 g29254 (.Q(n_74), 
	.B(B[9]), 
	.A(A[17]));
   EO2X3 g29255 (.Q(n_73), 
	.B(B[13]), 
	.A(A[19]));
   EO2X3 g29256 (.Q(n_72), 
	.B(B[3]), 
	.A(A[11]));
   EO2X3 g29257 (.Q(n_71), 
	.B(B[15]), 
	.A(A[20]));
   EO2X3 g29258 (.Q(n_70), 
	.B(B[15]), 
	.A(A[3]));
   EO2X3 g29259 (.Q(n_69), 
	.B(B[5]), 
	.A(A[12]));
   EO2X3 g29260 (.Q(n_68), 
	.B(B[5]), 
	.A(A[14]));
   EO2X3 g29261 (.Q(n_67), 
	.B(B[13]), 
	.A(A[10]));
   INX8 g29262 (.Q(n_65), 
	.A(n_66));
   EO2X3 g29263 (.Q(n_66), 
	.B(B[18]), 
	.A(B[17]));
   EO2X3 g29264 (.Q(n_64), 
	.B(B[9]), 
	.A(A[3]));
   EO2X3 g29265 (.Q(n_63), 
	.B(B[17]), 
	.A(A[17]));
   EO2X3 g29266 (.Q(n_62), 
	.B(B[17]), 
	.A(A[22]));
   EO2X3 g29267 (.Q(n_61), 
	.B(B[9]), 
	.A(A[5]));
   EN2X4 g29268 (.Q(n_60), 
	.B(B[11]), 
	.A(A[5]));
   EN2X4 g29269 (.Q(n_59), 
	.B(B[15]), 
	.A(A[17]));
   EO2X3 g29270 (.Q(n_58), 
	.B(B[5]), 
	.A(A[22]));
   EO2X3 g29271 (.Q(n_57), 
	.B(B[11]), 
	.A(A[6]));
   EN2X4 g29272 (.Q(n_56), 
	.B(B[21]), 
	.A(A[11]));
   EO2X3 g29273 (.Q(n_55), 
	.B(B[15]), 
	.A(A[11]));
   EO2X3 g29274 (.Q(n_54), 
	.B(B[7]), 
	.A(A[6]));
   EO2X3 g29275 (.Q(n_53), 
	.B(B[13]), 
	.A(A[3]));
   EO2X3 g29276 (.Q(n_52), 
	.B(B[17]), 
	.A(A[5]));
   EO2X3 g29277 (.Q(n_51), 
	.B(B[5]), 
	.A(A[9]));
   EO2X3 g29278 (.Q(n_50), 
	.B(B[7]), 
	.A(A[14]));
   INX4 g29279 (.Q(n_49), 
	.A(n_48));
   EN2X4 g29280 (.Q(n_48), 
	.B(B[19]), 
	.A(A[17]));
   EN2X4 g29281 (.Q(n_47), 
	.B(B[11]), 
	.A(A[23]));
   EN2X4 g29282 (.Q(n_46), 
	.B(B[3]), 
	.A(A[7]));
   EN2X4 g29283 (.Q(n_45), 
	.B(B[11]), 
	.A(A[21]));
   INX4 g29284 (.Q(n_44), 
	.A(n_43));
   EO2X3 g29285 (.Q(n_43), 
	.B(B[15]), 
	.A(A[15]));
   EO2X3 g29286 (.Q(n_42), 
	.B(B[13]), 
	.A(A[4]));
   EO2X3 g29287 (.Q(n_41), 
	.B(B[9]), 
	.A(A[1]));
   EO2X3 g29289 (.Q(n_40), 
	.B(B[9]), 
	.A(A[23]));
   EN2X4 g29290 (.Q(n_39), 
	.B(B[3]), 
	.A(A[5]));
   EO2X3 g29291 (.Q(n_38), 
	.B(B[13]), 
	.A(A[16]));
   INX4 g29292 (.Q(n_37), 
	.A(n_36));
   EO2X3 g29293 (.Q(n_36), 
	.B(B[17]), 
	.A(A[13]));
   EO2X3 g29294 (.Q(n_35), 
	.B(B[9]), 
	.A(A[16]));
   EN2X4 g29295 (.Q(n_34), 
	.B(B[7]), 
	.A(A[22]));
   EO2X3 g29296 (.Q(n_33), 
	.B(B[23]), 
	.A(A[13]));
   EO2X3 g29297 (.Q(n_32), 
	.B(B[23]), 
	.A(A[16]));
   EO2X3 g29298 (.Q(n_31), 
	.B(B[23]), 
	.A(A[10]));
   EO2X3 g29299 (.Q(n_30), 
	.B(B[23]), 
	.A(A[12]));
   EO2X3 g29300 (.Q(n_29), 
	.B(B[23]), 
	.A(A[15]));
   EO2X3 g29301 (.Q(n_28), 
	.B(B[23]), 
	.A(A[4]));
   EO2X3 g29302 (.Q(n_27), 
	.B(B[23]), 
	.A(A[1]));
   EO2X3 g29303 (.Q(n_26), 
	.B(B[23]), 
	.A(A[9]));
   NA2X4 g29306 (.Q(n_25), 
	.B(A[1]), 
	.A(B[23]));
   NA2X4 g29307 (.Q(n_24), 
	.B(A[16]), 
	.A(B[23]));
   NA2X4 g29308 (.Q(n_23), 
	.B(A[13]), 
	.A(B[23]));
   NA2X4 g29309 (.Q(n_22), 
	.B(A[15]), 
	.A(B[23]));
   NA2X4 g29310 (.Q(n_21), 
	.B(A[4]), 
	.A(B[23]));
   NA2X4 g29311 (.Q(n_20), 
	.B(A[10]), 
	.A(B[23]));
   NA2X4 g29312 (.Q(n_19), 
	.B(A[12]), 
	.A(B[23]));
   NA2X4 g29313 (.Q(n_18), 
	.B(A[9]), 
	.A(B[23]));
   INX8 g29315 (.Q(n_17), 
	.A(B[11]));
   INX8 g29316 (.Q(n_16), 
	.A(B[15]));
   INX8 g29317 (.Q(n_15), 
	.A(B[7]));
   INX8 g29321 (.Q(n_14), 
	.A(B[3]));
   INX8 g29322 (.Q(n_13), 
	.A(B[13]));
   EO2X3 g2 (.Q(n_12), 
	.B(n_1294), 
	.A(n_1288));
   EN2X4 g29326 (.Q(n_11), 
	.B(n_1282), 
	.A(n_1264));
   EO2X3 g29329 (.Q(n_10), 
	.B(n_1159), 
	.A(n_1081));
   EN2X4 g29332 (.Q(n_9), 
	.B(n_769), 
	.A(n_575));
   EN2X4 g29335 (.Q(n_8), 
	.B(n_777), 
	.A(n_743));
   EO2X3 g29338 (.Q(n_7), 
	.B(n_773), 
	.A(n_740));
   EO2X3 g29341 (.Q(n_6), 
	.B(n_782), 
	.A(n_746));
   EO2X3 g29344 (.Q(n_5), 
	.B(n_781), 
	.A(n_653));
   EO2X3 g29347 (.Q(n_4), 
	.B(n_783), 
	.A(n_528));
   EO2X2 g29350 (.Q(n_3), 
	.B(B[9]), 
	.A(B[10]));
   EO2X3 g29353 (.Q(n_2), 
	.B(B[21]), 
	.A(B[22]));
   AND2X4 g29356 (.Q(Z[0]), 
	.B(A[0]), 
	.A(B[0]));
   NO2I1X4 g29360 (.Q(n_0), 
	.B(B[0]), 
	.AN(B[1]));
endmodule

