#************************************************************************/
# Copyright        : (c) All Rights Reserved 
# Company          : X-FAB Semiconductor Foundries  
# Address          : Haarbergstr. 67,  D-99097 Erfurt, Germany 
#
# File             : xl035m3.lef 
# Description      : Layout Exchange Format
#                  
# Technology       : XL035M3
# Lib_version      : V 1.0.1
# Last Modified by : SKP
# DATE             : July 14, 2005 (r/c values corrected, tech.lef for FE) 
# 
#************************************************************************/
#  

VERSION 5.4 ;

NAMESCASESENSITIVE ON ;

BUSBITCHARS "[]" ;

UNITS
    DATABASE MICRONS 1000  ;
	RESISTANCE OHMS 10 ;
	ARTEMKA MOLODEC 5 ;	
END UNITS

MANUFACTURINGGRID 0.025 ;

LAYER M1M
    TYPE ROUTING ;
    WIDTH 0.5 ;
    SPACING 0.45 ;
    PITCH 1.3 ;
    DIRECTION HORIZONTAL ;
    CAPACITANCE CPERSQDIST 0.0000400000 ;
    RESISTANCE RPERSQ 0.12000000 ;
    EDGECAPACITANCE 0.0000460000 ;
    ANTENNAAREARATIO 100 ;
    ANTENNADIFFAREARATIO 9999999 ; 
END M1M

LAYER V1M
    TYPE CUT ;
END V1M
 
LAYER M2M
    TYPE ROUTING ;
    WIDTH 0.6 ;
    SPACING 0.5 ;
    PITCH 1.4 ;
    DIRECTION VERTICAL ;
    CAPACITANCE CPERSQDIST 0.0000134000 ;
    RESISTANCE RPERSQ 0.12000000 ;
    EDGECAPACITANCE 0.0000300000 ;
    ANTENNAAREARATIO 100 ;
    ANTENNADIFFAREARATIO 9999999 ; 
END M2M
 
LAYER V2M
    TYPE CUT ;
END V2M
 
LAYER M3M
    TYPE ROUTING ;
    WIDTH 0.6 ;
    SPACING 0.6 ;
    PITCH 1.3 ;
    DIRECTION HORIZONTAL ;
    CAPACITANCE CPERSQDIST 0.0000086000 ;
    RESISTANCE RPERSQ 0.12000000 ;
    EDGECAPACITANCE 0.0000240000 ;
    ANTENNAAREARATIO 100 ;
    ANTENNADIFFAREARATIO 9999999 ; 
END M3M

# Via Met1-Met2 for normal routing
VIA CLVIA1 DEFAULT
    RESISTANCE 6 ;
    FOREIGN CLVIA1 ;
    LAYER M1M ;
        RECT -0.450000 -0.450000 0.450000 0.450000 ;
    LAYER V1M ;
        RECT -0.250000 -0.250000 0.250000 0.250000 ;
    LAYER M2M ;
        RECT -0.400000 -0.400000 0.400000 0.400000 ;
END CLVIA1

# Via Met2-Met3 for normal routing
VIA CLVIA2 DEFAULT
    RESISTANCE 6 ;
    FOREIGN CLVIA2 ;
    LAYER M2M ;
        RECT -0.450000 -0.450000 0.450000 0.450000 ;
    LAYER V2M ;
        RECT -0.250000 -0.250000 0.250000 0.250000 ;
    LAYER M3M ;
        RECT -0.400000 -0.400000 0.400000 0.400000 ;
END CLVIA2

# Rule Via (needed for DEF import to DFII)
VIA ruleV1
        LAYER M1M ;
          RECT -0.950000 -0.450000 0.950000 0.450000 ;
        LAYER V1M ;
          RECT -0.750000 -0.250000 -0.250000 0.250000 ;
          RECT 0.250000 -0.250000 0.750000 0.250000 ;
        LAYER M2M ;
          RECT -0.900000 -0.400000 0.900000 0.400000 ;
END ruleV1

# Rule Via (needed for DEF import to DFII)
VIA ruleV2
        LAYER M2M ;
          RECT -0.950000 -0.450000 0.950000 0.450000 ;
        LAYER V2M ;
          RECT -0.750000 -0.250000 -0.250000 0.250000 ;
          RECT 0.250000 -0.250000 0.750000 0.250000 ;
        LAYER M3M ;
          RECT -0.900000 -0.400000 0.900000 0.400000 ;
END ruleV2

# V1 Array for Wide-Met1/Wide-Met2
VIARULE V1M12W GENERATE
    LAYER M2M ;
       DIRECTION VERTICAL ; 
       WIDTH 10 TO 1000.0 ; 
       OVERHANG 0.15 ;
       METALOVERHANG 0.00 ;
       ENCLOSURE 1 2;

    LAYER M1M ;
        DIRECTION HORIZONTAL ; 
        WIDTH 10 TO 1000.0 ; 
        OVERHANG 0.15 ;
        METALOVERHANG 0.05 ;
	ENCLOSURE 3 4;

    LAYER V1M ;
        RECT -0.250000 -0.250000 0.250000 0.250000 ;
        SPACING 0.950000 BY 0.950000 ;
    RESISTANCE 6 ;
END V1M12W

# V1 Array for Wide-Met1/Met2
# normal routing direction Met1 horizontal/Met2 vertical 
VIARULE V1WM1M2 GENERATE
    LAYER M2M ;
        DIRECTION VERTICAL ; 
        OVERHANG 0.15 ;
        METALOVERHANG 0.00 ;

    LAYER M1M ;
        DIRECTION HORIZONTAL ; 
        WIDTH 10 TO 1000.0 ; 
        OVERHANG 0.15 ;
        METALOVERHANG 0.05 ;

    LAYER V1M ;
        RECT -0.250000 -0.250000 0.250000 0.250000 ;
        SPACING 0.950000 BY 0.950000 ;
    RESISTANCE 6 ;
END V1WM1M2

# V1 Array for Met1/Wide-Met2
# Normal routing direction Met1 horizontal / Met2 vertical
VIARULE V1M1WM2 GENERATE
    LAYER M2M ;
        DIRECTION VERTICAL ; 
        WIDTH 10 TO 1000.0 ; 
        OVERHANG 0.15 ;
        METALOVERHANG 0.00 ;

    LAYER M1M ;
        DIRECTION HORIZONTAL ; 
        OVERHANG 0.15 ;
        METALOVERHANG 0.05 ;

    LAYER V1M ;
        RECT -0.250000 -0.250000 0.250000 0.250000 ;
        SPACING 0.950000 BY 0.950000 ;
    RESISTANCE 6 ;
END V1M1WM2

# V2 Array for Wide-Met2/Wide-Met3
VIARULE V2M23W GENERATE
    LAYER M3M ;
       DIRECTION VERTICAL ; 
       WIDTH 10 TO 1000.0 ; 
       OVERHANG 0.15 ;
       METALOVERHANG 0.00 ;

    LAYER M2M ;
        DIRECTION HORIZONTAL ; 
        WIDTH 10 TO 1000.0 ; 
        OVERHANG 0.15 ;
        METALOVERHANG 0.05 ;

    LAYER V2M ;
        RECT -0.250000 -0.250000 0.250000 0.250000 ;
        SPACING 0.950000 BY 0.950000 ;
    RESISTANCE 6 ;
END V2M23W

# V2 Array for Wide-Met2/Met3
# normal routing direction Met2 horizontal/Met3 vertical 
VIARULE V2WM2M3 GENERATE
    LAYER M3M ;
        DIRECTION VERTICAL ; 
        OVERHANG 0.15 ;
        METALOVERHANG 0.00 ;

    LAYER M2M ;
        DIRECTION HORIZONTAL ; 
        WIDTH 10 TO 1000.0 ; 
        OVERHANG 0.15 ;
        METALOVERHANG 0.05 ;

    LAYER V2M ;
        RECT -0.250000 -0.250000 0.250000 0.250000 ;
        SPACING 0.950000 BY 0.950000 ;
    RESISTANCE 6 ;
END V2WM2M3

# V2 Array for Met2/Wide-Met3
# Normal routing direction Met2 horizontal / Met3 vertical
VIARULE V2M2WM3 GENERATE
    LAYER M3M ;
        DIRECTION VERTICAL ; 
        WIDTH 10 TO 1000.0 ; 
        OVERHANG 0.15 ;
        METALOVERHANG 0.00 ;

    LAYER M2M ;
        DIRECTION HORIZONTAL ; 
        OVERHANG 0.15 ;
        METALOVERHANG 0.05 ;

    LAYER V2M ;
        RECT -0.250000 -0.250000 0.250000 0.250000 ;
        SPACING 0.950000 BY 0.950000 ;
    RESISTANCE 6 ;
END V2M2WM3
 

# V1 Array for Met1/Met2
VIARULE V1M12 GENERATE
    LAYER M2M ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.15 ;
        METALOVERHANG 0.00 ;

    LAYER M1M ;
        DIRECTION VERTICAL ;
        OVERHANG 0.15 ;
        METALOVERHANG 0.05 ;

    LAYER V1M ;
        RECT -0.250000 -0.250000 0.250000 0.250000 ;
        SPACING 0.950000 BY 0.950000 ;
    RESISTANCE 6 ;
END V1M12

# V2 Array for Met2/Met3
VIARULE V2M23 GENERATE
    LAYER M3M ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.15 ;
        METALOVERHANG 0.00 ;

    LAYER M2M ;
        DIRECTION VERTICAL ;
        OVERHANG 0.15 ;
        METALOVERHANG 0.05 ;

    LAYER V2M ;
        RECT -0.250000 -0.250000 0.250000 0.250000 ;
        SPACING 0.950000 BY 0.950000 ;
    RESISTANCE 6 ;
END V2M23

# Turn Vias
VIARULE TURN1 GENERATE
    LAYER M1M ;
        DIRECTION vertical ;
 
    LAYER M1M ;
        DIRECTION horizontal ;
END TURN1
 
VIARULE TURN2 GENERATE
    LAYER M2M ;
        DIRECTION vertical ;
 
    LAYER M2M ;
        DIRECTION horizontal ;
END TURN2
 
VIARULE TURN3 GENERATE
    LAYER M3M ;
        DIRECTION vertical ;
 
    LAYER M3M ;
        DIRECTION horizontal ;
END TURN3
 
 
SPACING
    SAMENET M1M M1M 0.45 STACK ;
    SAMENET M2M M2M 0.50 STACK ;
    SAMENET M3M M3M 0.50 STACK ;
    SAMENET V1M V1M 0.45 STACK ;
    SAMENET V2M V2M 0.45 STACK ;
END SPACING
  
END LIBRARY
