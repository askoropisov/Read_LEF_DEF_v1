#$Id: mksoi018std9t1v8.lef 1427 2020-11-24 13:59:11Z silin $
#******
# Preview export LEF
#
#	 Preview sub-version 5.10.41.500.6.151
#
# REF LIBS: mksoi018std9t1v8
# TECH LIB NAME: LibMikron_SOI_018_6M
# TECH FILE NAME: techfile.cds
#******

VERSION 5.7 ;

DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

UNITS
    DATABASE MICRONS 100  ;
END UNITS

 MANUFACTURINGGRID    0.010000 ;
SITE CORE
    SYMMETRY X Y  ;
    CLASS CORE  ;
    SIZE 0.64 BY 5.76 ;
END CORE

MACRO tinvh_8
    CLASS CORE ;
    FOREIGN tinvh_8 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.24 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.72 ;
        END
    END a
    PIN en
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.06  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 1.76 2.72 ;
        END
    END en
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.74  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  5.84 1.54 5.72 1.54 5.60 1.66 5.60 3.90 3.64 3.90 3.64 3.58
                 5.28 3.58 5.28 1.46 5.52 1.22 5.84 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  10.24 0.90 9.36 0.90 9.36 1.14 9.04 1.14 9.04 0.90 8.64 0.90
                 8.64 1.14 8.32 1.14 8.32 0.90 7.22 0.90 7.22 1.14 6.90 1.14
                 6.90 0.90 6.54 0.90 6.54 1.14 6.22 1.14 6.22 0.90 5.14 0.90
                 5.14 1.14 4.82 1.14 4.82 0.90 1.28 0.90 1.28 1.58 0.96 1.58
                 0.96 0.90 0.00 0.90 0.00 -0.90 10.24 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 10.24 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  10.06 4.10 9.74 4.10 9.74 1.78 8.56 1.78 8.56 2.65 7.46 2.65
                 7.46 2.33 8.24 2.33 8.24 1.46 9.74 1.46 9.74 1.22 10.06 1.22 ;
        POLYGON  9.27 4.54 0.16 4.54 0.16 1.26 0.50 1.26 0.50 1.58 0.48 1.58
                 0.48 3.10 1.94 3.10 1.94 3.42 0.48 3.42 0.48 4.22 8.95 4.22
                 8.95 2.66 8.88 2.66 8.88 2.34 9.27 2.34 ;
        RECT  7.42 3.58 8.42 3.90 ;
        POLYGON  7.92 1.78 7.14 1.78 7.14 2.34 7.04 2.34 7.04 3.90 6.72 3.90
                 6.72 2.98 5.93 2.98 5.93 2.66 6.72 2.66 6.72 2.02 6.82 2.02
                 6.82 1.46 7.92 1.46 ;
        POLYGON  4.46 2.89 2.58 2.89 2.58 3.90 2.26 3.90 2.26 2.57 3.20 2.57
                 3.20 1.22 3.52 1.22 3.52 2.57 4.46 2.57 ;
        RECT  1.82 1.22 2.84 1.54 ;
    END
END tinvh_8

MACRO tinvh_64
    CLASS CORE ;
    FOREIGN tinvh_64 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 32.64 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.33 1.12 3.04 ;
        END
    END a
    PIN en
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.08 2.62 9.25 2.62 9.25 2.30 9.76 2.30 9.76 2.08 10.08 2.08 ;
        END
    END en
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 16.39  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  22.34 3.90 19.11 3.90 19.11 1.78 16.76 1.78 16.76 3.58
                 19.11 3.58 19.11 3.90 16.44 3.90 16.44 1.78 13.92 1.78
                 13.92 3.58 16.44 3.58 16.44 3.90 13.60 3.90 13.60 1.78
                 11.16 1.78 11.16 3.58 13.60 3.58 13.60 3.90 9.37 3.90
                 9.37 3.58 10.84 3.58 10.84 1.46 20.96 1.46 20.96 1.78
                 19.43 1.78 19.43 3.58 22.34 3.58 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  32.64 0.90 31.37 0.90 31.37 1.16 31.05 1.16 31.05 0.90
                 28.95 0.90 28.95 1.16 28.63 1.16 28.63 0.90 27.55 0.90
                 27.55 1.16 27.23 1.16 27.23 0.90 26.15 0.90 26.15 1.16
                 25.83 1.16 25.83 0.90 24.75 0.90 24.75 1.16 24.43 1.16
                 24.43 0.90 21.66 0.90 21.66 1.14 21.34 1.14 21.34 0.90
                 20.26 0.90 20.26 1.14 19.94 1.14 19.94 0.90 18.86 0.90
                 18.86 1.14 18.54 1.14 18.54 0.90 17.46 0.90 17.46 1.14
                 17.14 1.14 17.14 0.90 16.06 0.90 16.06 1.14 15.74 1.14
                 15.74 0.90 14.66 0.90 14.66 1.14 14.34 1.14 14.34 0.90
                 13.26 0.90 13.26 1.14 12.94 1.14 12.94 0.90 11.86 0.90
                 11.86 1.14 11.54 1.14 11.54 0.90 10.46 0.90 10.46 1.14
                 10.14 1.14 10.14 0.90 1.20 0.90 1.20 1.32 0.88 1.32 0.88 0.90
                 0.00 0.90 0.00 -0.90 32.64 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 32.64 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  32.07 1.80 30.67 1.80 30.67 3.43 32.07 3.43 32.07 4.54
                 31.75 4.54 31.75 3.75 30.67 3.75 30.67 4.54 30.35 4.54
                 30.35 2.62 28.33 2.62 28.33 2.30 30.35 2.30 30.35 1.48
                 32.07 1.48 ;
        POLYGON  29.99 3.85 29.67 3.85 29.67 3.26 28.59 3.26 28.59 3.85
                 28.27 3.85 28.27 3.26 27.19 3.26 27.19 3.85 26.87 3.85
                 26.87 1.92 23.25 1.92 23.25 2.81 20.26 2.81 20.26 2.48
                 22.93 2.48 22.93 1.60 29.65 1.60 29.65 1.92 27.19 1.92
                 27.19 2.94 29.99 2.94 ;
        RECT  23.39 4.17 29.33 4.49 ;
        POLYGON  24.77 2.60 24.14 2.60 24.14 3.67 23.07 3.67 23.07 4.53
                 23.00 4.53 23.00 4.54 0.18 4.54 0.18 3.26 0.50 3.26 0.50 4.22
                 1.58 4.22 1.58 1.96 0.18 1.96 0.18 1.64 1.90 1.64 1.90 2.90
                 2.98 2.90 2.98 3.22 1.90 3.22 1.90 4.22 22.75 4.22 22.75 3.35
                 23.82 3.35 23.82 2.28 24.77 2.28 ;
        POLYGON  10.32 3.26 8.18 3.26 8.18 3.90 2.26 3.90 2.26 3.58 7.86 3.58
                 7.86 2.34 5.74 2.34 5.74 2.02 8.54 2.02 8.54 1.34 8.86 1.34
                 8.86 2.34 8.18 2.34 8.18 2.94 10.32 2.94 ;
        RECT  2.26 1.32 8.16 1.64 ;
    END
END tinvh_64

MACRO tinvh_6
    CLASS CORE ;
    FOREIGN tinvh_6 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.24 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.72 ;
        END
    END a
    PIN en
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.06  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 1.76 2.72 ;
        END
    END en
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.62  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  5.84 1.54 5.72 1.54 5.60 1.66 5.60 3.90 3.64 3.90 3.64 3.58
                 5.28 3.58 5.28 1.46 5.52 1.22 5.84 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  10.24 0.90 9.36 0.90 9.36 1.14 9.04 1.14 9.04 0.90 8.64 0.90
                 8.64 1.14 8.32 1.14 8.32 0.90 7.22 0.90 7.22 1.14 6.90 1.14
                 6.90 0.90 6.54 0.90 6.54 1.14 6.22 1.14 6.22 0.90 5.14 0.90
                 5.14 1.14 4.82 1.14 4.82 0.90 1.28 0.90 1.28 1.58 0.96 1.58
                 0.96 0.90 0.00 0.90 0.00 -0.90 10.24 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 10.24 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  10.06 4.10 9.74 4.10 9.74 1.78 8.56 1.78 8.56 2.65 7.46 2.65
                 7.46 2.33 8.24 2.33 8.24 1.46 9.74 1.46 9.74 1.22 10.06 1.22 ;
        POLYGON  9.27 4.54 0.16 4.54 0.16 1.26 0.50 1.26 0.50 1.58 0.48 1.58
                 0.48 3.10 1.94 3.10 1.94 3.42 0.48 3.42 0.48 4.22 8.95 4.22
                 8.95 2.66 8.88 2.66 8.88 2.34 9.27 2.34 ;
        RECT  7.42 3.58 8.42 3.90 ;
        POLYGON  7.92 1.78 7.14 1.78 7.14 2.34 7.04 2.34 7.04 3.90 6.72 3.90
                 6.72 2.98 5.93 2.98 5.93 2.66 6.72 2.66 6.72 2.02 6.82 2.02
                 6.82 1.46 7.92 1.46 ;
        POLYGON  4.46 2.89 2.58 2.89 2.58 3.90 2.26 3.90 2.26 2.57 3.20 2.57
                 3.20 1.22 3.52 1.22 3.52 2.57 4.46 2.57 ;
        RECT  1.82 1.22 2.84 1.54 ;
    END
END tinvh_6

MACRO tinvh_48
    CLASS CORE ;
    FOREIGN tinvh_48 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 31.36 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  0.80 2.66 0.16 2.66 0.16 2.08 0.48 2.08 0.48 2.34 0.80 2.34 ;
        END
    END a
    PIN en
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.97  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.44 2.62 8.79 2.62 8.79 2.30 9.12 2.30 9.12 2.08 9.44 2.08 ;
        END
    END en
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 15.82  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  21.88 3.90 18.65 3.90 18.65 1.78 16.30 1.78 16.30 3.58
                 18.65 3.58 18.65 3.90 15.98 3.90 15.98 1.78 13.28 1.78
                 13.28 3.58 15.98 3.58 15.98 3.90 12.96 3.90 12.96 1.78
                 10.70 1.78 10.70 3.58 12.96 3.58 12.96 3.90 8.91 3.90
                 8.91 3.58 10.38 3.58 10.38 1.46 20.50 1.46 20.50 1.78
                 18.97 1.78 18.97 3.58 21.88 3.58 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  31.36 0.90 30.21 0.90 30.21 1.16 29.89 1.16 29.89 0.90
                 28.49 0.90 28.49 1.16 28.17 1.16 28.17 0.90 27.09 0.90
                 27.09 1.16 26.77 1.16 26.77 0.90 25.69 0.90 25.69 1.16
                 25.37 1.16 25.37 0.90 24.29 0.90 24.29 1.16 23.97 1.16
                 23.97 0.90 21.20 0.90 21.20 1.14 20.88 1.14 20.88 0.90
                 19.80 0.90 19.80 1.14 19.48 1.14 19.48 0.90 18.40 0.90
                 18.40 1.14 18.08 1.14 18.08 0.90 17.00 0.90 17.00 1.14
                 16.68 1.14 16.68 0.90 15.60 0.90 15.60 1.14 15.28 1.14
                 15.28 0.90 14.20 0.90 14.20 1.14 13.88 1.14 13.88 0.90
                 12.80 0.90 12.80 1.14 12.48 1.14 12.48 0.90 11.40 0.90
                 11.40 1.14 11.08 1.14 11.08 0.90 10.00 0.90 10.00 1.14
                 9.68 1.14 9.68 0.90 0.74 0.90 0.74 1.32 0.42 1.32 0.42 0.90
                 0.00 0.90 0.00 -0.90 31.36 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 31.36 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  30.91 4.54 30.59 4.54 30.59 2.62 27.87 2.62 27.87 2.30
                 30.59 2.30 30.59 1.48 30.91 1.48 ;
        POLYGON  29.53 3.85 29.21 3.85 29.21 3.26 28.13 3.26 28.13 3.85
                 27.81 3.85 27.81 3.26 26.73 3.26 26.73 3.85 26.41 3.85
                 26.41 1.92 22.79 1.92 22.79 2.81 19.80 2.81 19.80 2.48
                 22.47 2.48 22.47 1.60 29.19 1.60 29.19 1.92 26.73 1.92
                 26.73 2.94 29.53 2.94 ;
        RECT  22.93 4.17 28.87 4.49 ;
        POLYGON  24.31 2.60 23.68 2.60 23.68 3.67 22.61 3.67 22.61 4.53
                 22.54 4.53 22.54 4.54 0.47 4.54 0.47 4.22 1.12 4.22 1.12 1.64
                 1.44 1.64 1.44 2.90 2.52 2.90 2.52 3.22 1.44 3.22 1.44 4.22
                 22.29 4.22 22.29 3.35 23.36 3.35 23.36 2.28 24.31 2.28 ;
        POLYGON  9.86 3.26 7.72 3.26 7.72 3.90 1.80 3.90 1.80 3.58 7.40 3.58
                 7.40 2.34 5.28 2.34 5.28 2.02 8.08 2.02 8.08 1.34 8.40 1.34
                 8.40 2.34 7.72 2.34 7.72 2.94 9.86 2.94 ;
        RECT  1.80 1.32 7.70 1.64 ;
    END
END tinvh_48

MACRO tinvh_4
    CLASS CORE ;
    FOREIGN tinvh_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.96 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.72 ;
        END
    END a
    PIN en
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.06  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 1.76 2.72 ;
        END
    END en
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.64  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  5.19 1.54 5.07 1.54 4.98 1.63 4.98 3.90 4.39 3.90 4.39 3.58
                 4.66 3.58 4.66 2.40 4.64 2.40 4.64 2.08 4.66 2.08 4.66 1.43
                 4.87 1.22 5.19 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.96 0.90 8.08 0.90 8.08 1.14 7.76 1.14 7.76 0.90 7.36 0.90
                 7.36 1.14 7.04 1.14 7.04 0.90 5.87 0.90 5.87 1.14 5.55 1.14
                 5.55 0.90 4.49 0.90 4.49 1.14 4.17 1.14 4.17 0.90 1.28 0.90
                 1.28 1.58 0.96 1.58 0.96 0.90 0.00 0.90 0.00 -0.90 8.96 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 8.96 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  8.78 4.10 8.46 4.10 8.46 1.78 7.21 1.78 7.21 2.65 6.18 2.65
                 6.18 2.33 6.89 2.33 6.89 1.46 8.46 1.46 8.46 1.22 8.78 1.22 ;
        POLYGON  7.99 4.54 0.16 4.54 0.16 1.26 0.50 1.26 0.50 1.58 0.48 1.58
                 0.48 3.10 1.94 3.10 1.94 3.42 0.48 3.42 0.48 4.22 7.67 4.22
                 7.67 2.66 7.56 2.66 7.56 2.34 7.99 2.34 ;
        RECT  6.14 3.58 7.14 3.90 ;
        POLYGON  6.57 1.78 5.86 1.78 5.86 2.34 5.76 2.34 5.76 3.90 5.44 3.90
                 5.44 2.34 5.30 2.34 5.30 2.02 5.54 2.02 5.54 1.46 6.57 1.46 ;
        POLYGON  4.34 2.96 2.58 2.96 2.58 3.90 2.26 3.90 2.26 2.64 3.20 2.64
                 3.20 1.22 3.52 1.22 3.52 2.64 4.34 2.64 ;
        RECT  1.82 1.22 2.84 1.54 ;
    END
END tinvh_4

MACRO tinvh_32
    CLASS CORE ;
    FOREIGN tinvh_32 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 17.92 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.86 1.12 2.50 ;
        END
    END a
    PIN en
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.83  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 1.86 1.78 2.48 ;
        END
    END en
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 8.89  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.36 3.90 9.77 3.90 9.77 1.78 7.52 1.78 7.52 3.58 9.77 3.58
                 9.77 3.90 5.04 3.90 5.04 3.58 7.20 3.58 7.20 1.78 6.62 1.78
                 6.62 1.46 11.14 1.46 11.14 1.78 10.09 1.78 10.09 3.58
                 12.36 3.58 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  17.92 0.90 15.46 0.90 15.46 1.14 15.14 1.14 15.14 0.90
                 14.06 0.90 14.06 1.14 13.74 1.14 13.74 0.90 11.84 0.90
                 11.84 1.14 11.52 1.14 11.52 0.90 10.44 0.90 10.44 1.14
                 10.12 1.14 10.12 0.90 9.04 0.90 9.04 1.14 8.72 1.14 8.72 0.90
                 7.64 0.90 7.64 1.14 7.32 1.14 7.32 0.90 6.24 0.90 6.24 1.14
                 5.92 1.14 5.92 0.90 1.32 0.90 1.32 1.54 1.00 1.54 1.00 0.90
                 0.00 0.90 0.00 -0.90 17.92 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 17.92 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  17.70 4.10 17.38 4.10 17.38 2.62 14.10 2.62 14.10 2.30
                 17.38 2.30 17.38 1.22 17.70 1.22 ;
        POLYGON  16.91 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 2.94 1.88 2.94 1.88 3.26 0.48 3.26 0.48 4.22 16.59 4.22
                 16.59 3.26 14.56 3.26 14.56 2.94 16.91 2.94 ;
        POLYGON  16.16 1.78 13.76 1.78 13.76 3.26 13.42 3.26 13.42 2.80
                 10.54 2.80 10.54 2.48 13.42 2.48 13.42 1.78 13.04 1.78
                 13.04 1.46 16.16 1.46 ;
        RECT  12.72 3.58 16.02 3.90 ;
        POLYGON  6.76 3.26 4.68 3.26 4.68 3.90 4.36 3.90 4.36 3.26 3.28 3.26
                 3.28 3.90 1.56 3.90 1.56 3.58 2.96 3.58 2.96 2.94 3.90 2.94
                 3.90 1.86 4.22 1.86 4.22 2.94 6.76 2.94 ;
        RECT  1.82 1.22 4.92 1.54 ;
    END
END tinvh_32

MACRO tinvh_3
    CLASS CORE ;
    FOREIGN tinvh_3 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.96 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.45  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.72 ;
        END
    END a
    PIN en
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.02  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 1.76 2.72 ;
        END
    END en
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.58  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  5.19 1.54 5.07 1.54 4.98 1.63 4.98 3.90 4.39 3.90 4.39 3.58
                 4.66 3.58 4.66 2.40 4.64 2.40 4.64 2.08 4.66 2.08 4.66 1.43
                 4.87 1.22 5.19 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.96 0.90 8.08 0.90 8.08 1.14 7.76 1.14 7.76 0.90 7.36 0.90
                 7.36 1.14 7.04 1.14 7.04 0.90 5.87 0.90 5.87 1.14 5.55 1.14
                 5.55 0.90 4.49 0.90 4.49 1.14 4.17 1.14 4.17 0.90 1.28 0.90
                 1.28 1.58 0.96 1.58 0.96 0.90 0.00 0.90 0.00 -0.90 8.96 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 8.96 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  8.78 4.34 8.46 4.34 8.46 1.78 7.21 1.78 7.21 2.65 6.18 2.65
                 6.18 2.33 6.89 2.33 6.89 1.46 8.46 1.46 8.46 1.22 8.78 1.22 ;
        POLYGON  7.99 4.54 0.16 4.54 0.16 1.26 0.50 1.26 0.50 1.58 0.48 1.58
                 0.48 3.10 1.94 3.10 1.94 3.42 0.48 3.42 0.48 4.22 7.67 4.22
                 7.67 2.66 7.56 2.66 7.56 2.34 7.99 2.34 ;
        RECT  6.14 3.58 7.14 3.90 ;
        POLYGON  6.57 1.78 5.86 1.78 5.86 2.34 5.76 2.34 5.76 3.90 5.44 3.90
                 5.44 2.34 5.30 2.34 5.30 2.02 5.54 2.02 5.54 1.46 6.57 1.46 ;
        POLYGON  4.34 2.96 2.58 2.96 2.58 3.90 2.26 3.90 2.26 2.64 3.20 2.64
                 3.20 1.22 3.52 1.22 3.52 2.64 4.34 2.64 ;
        RECT  1.82 1.22 2.84 1.54 ;
    END
END tinvh_3

MACRO tinvh_24
    CLASS CORE ;
    FOREIGN tinvh_24 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 17.92 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.86 1.12 2.50 ;
        END
    END a
    PIN en
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.83  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 1.86 1.78 2.48 ;
        END
    END en
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 8.56  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.36 3.90 9.77 3.90 9.77 1.78 7.52 1.78 7.52 3.58 9.77 3.58
                 9.77 3.90 5.04 3.90 5.04 3.58 7.20 3.58 7.20 1.78 6.62 1.78
                 6.62 1.46 11.14 1.46 11.14 1.78 10.09 1.78 10.09 3.58
                 12.36 3.58 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  17.92 0.90 15.46 0.90 15.46 1.14 15.14 1.14 15.14 0.90
                 14.06 0.90 14.06 1.14 13.74 1.14 13.74 0.90 11.84 0.90
                 11.84 1.14 11.52 1.14 11.52 0.90 10.44 0.90 10.44 1.14
                 10.12 1.14 10.12 0.90 9.04 0.90 9.04 1.14 8.72 1.14 8.72 0.90
                 7.64 0.90 7.64 1.14 7.32 1.14 7.32 0.90 6.24 0.90 6.24 1.14
                 5.92 1.14 5.92 0.90 1.32 0.90 1.32 1.54 1.00 1.54 1.00 0.90
                 0.00 0.90 0.00 -0.90 17.92 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 17.92 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  17.70 4.10 17.38 4.10 17.38 2.62 14.10 2.62 14.10 2.30
                 17.38 2.30 17.38 1.22 17.70 1.22 ;
        POLYGON  16.91 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 2.94 1.88 2.94 1.88 3.26 0.48 3.26 0.48 4.22 16.59 4.22
                 16.59 3.26 14.56 3.26 14.56 2.94 16.91 2.94 ;
        POLYGON  16.16 1.78 13.76 1.78 13.76 3.26 13.42 3.26 13.42 2.80
                 10.54 2.80 10.54 2.48 13.42 2.48 13.42 1.78 13.04 1.78
                 13.04 1.46 16.16 1.46 ;
        RECT  12.72 3.58 16.02 3.90 ;
        POLYGON  6.76 3.26 4.68 3.26 4.68 3.90 4.36 3.90 4.36 3.26 3.28 3.26
                 3.28 3.90 1.56 3.90 1.56 3.58 2.96 3.58 2.96 2.94 3.90 2.94
                 3.90 1.86 4.22 1.86 4.22 2.94 6.76 2.94 ;
        RECT  1.82 1.22 4.92 1.54 ;
    END
END tinvh_24

MACRO tinvh_20
    CLASS CORE ;
    FOREIGN tinvh_20 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.64 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.86 1.12 2.50 ;
        END
    END a
    PIN en
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 1.86 1.78 2.48 ;
        END
    END en
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 7.22  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.96 3.90 8.90 3.90 8.90 1.78 7.52 1.78 7.52 3.58 8.90 3.58
                 8.90 3.90 5.04 3.90 5.04 3.58 7.20 3.58 7.20 1.78 6.08 1.78
                 6.08 1.46 10.60 1.46 10.60 1.78 9.22 1.78 9.22 3.58 10.96 3.58 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 0.90 14.18 0.90 14.18 1.14 13.86 1.14 13.86 0.90
                 12.78 0.90 12.78 1.14 12.46 1.14 12.46 0.90 11.30 0.90
                 11.30 1.14 10.98 1.14 10.98 0.90 9.90 0.90 9.90 1.14 9.58 1.14
                 9.58 0.90 8.50 0.90 8.50 1.14 8.18 1.14 8.18 0.90 7.10 0.90
                 7.10 1.14 6.78 1.14 6.78 0.90 5.70 0.90 5.70 1.14 5.38 1.14
                 5.38 0.90 0.00 0.90 0.00 -0.90 16.64 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 16.64 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  16.42 4.39 16.10 4.39 16.10 2.62 12.82 2.62 12.82 2.30
                 16.10 2.30 16.10 1.22 16.42 1.22 ;
        POLYGON  15.63 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 2.94 1.88 2.94 1.88 3.26 0.48 3.26 0.48 4.22 15.31 4.22
                 15.31 3.26 13.28 3.26 13.28 2.94 15.63 2.94 ;
        POLYGON  14.88 1.78 12.48 1.78 12.48 3.26 12.14 3.26 12.14 2.80
                 10.00 2.80 10.00 2.48 12.14 2.48 12.14 1.78 11.76 1.78
                 11.76 1.46 14.88 1.46 ;
        RECT  11.44 3.58 14.74 3.90 ;
        POLYGON  6.77 3.26 4.68 3.26 4.68 3.90 4.36 3.90 4.36 3.26 3.28 3.26
                 3.28 3.90 1.56 3.90 1.56 3.58 2.96 3.58 2.96 2.94 3.90 2.94
                 3.90 1.86 4.22 1.86 4.22 2.94 6.77 2.94 ;
        RECT  1.82 1.22 4.92 1.54 ;
    END
END tinvh_20

MACRO tinvh_2
    CLASS CORE ;
    FOREIGN tinvh_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.96 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.45  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.72 ;
        END
    END a
    PIN en
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.02  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 1.76 2.72 ;
        END
    END en
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.38  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  5.19 1.54 5.07 1.54 4.98 1.63 4.98 3.90 4.39 3.90 4.39 3.58
                 4.66 3.58 4.66 2.40 4.64 2.40 4.64 2.08 4.66 2.08 4.66 1.43
                 4.87 1.22 5.19 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.96 0.90 8.08 0.90 8.08 1.14 7.76 1.14 7.76 0.90 7.36 0.90
                 7.36 1.14 7.04 1.14 7.04 0.90 5.87 0.90 5.87 1.14 5.55 1.14
                 5.55 0.90 4.49 0.90 4.49 1.14 4.17 1.14 4.17 0.90 1.28 0.90
                 1.28 1.58 0.96 1.58 0.96 0.90 0.00 0.90 0.00 -0.90 8.96 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 8.96 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  8.78 4.34 8.46 4.34 8.46 1.78 7.21 1.78 7.21 2.65 6.18 2.65
                 6.18 2.33 6.89 2.33 6.89 1.46 8.46 1.46 8.46 1.22 8.78 1.22 ;
        POLYGON  7.99 4.54 0.16 4.54 0.16 1.26 0.50 1.26 0.50 1.58 0.48 1.58
                 0.48 3.10 1.94 3.10 1.94 3.42 0.48 3.42 0.48 4.22 7.67 4.22
                 7.67 2.66 7.56 2.66 7.56 2.34 7.99 2.34 ;
        RECT  6.14 3.58 7.14 3.90 ;
        POLYGON  6.57 1.78 5.86 1.78 5.86 2.34 5.76 2.34 5.76 3.90 5.44 3.90
                 5.44 2.34 5.30 2.34 5.30 2.02 5.54 2.02 5.54 1.46 6.57 1.46 ;
        POLYGON  4.34 2.96 2.58 2.96 2.58 3.90 2.26 3.90 2.26 2.64 3.20 2.64
                 3.20 1.22 3.52 1.22 3.52 2.64 4.34 2.64 ;
        RECT  1.82 1.22 2.84 1.54 ;
    END
END tinvh_2

MACRO tinvh_16
    CLASS CORE ;
    FOREIGN tinvh_16 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.52 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.72 ;
        END
    END a
    PIN en
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.06  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 1.76 2.72 ;
        END
    END en
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.44  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  6.94 1.78 5.60 1.78 5.60 3.58 6.78 3.58 6.78 3.90 3.64 3.90
                 3.64 3.58 5.28 3.58 5.28 1.78 5.22 1.78 5.22 1.46 6.94 1.46 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  11.52 0.90 10.46 0.90 10.46 1.14 10.14 1.14 10.14 0.90
                 9.74 0.90 9.74 1.14 9.42 1.14 9.42 0.90 8.32 0.90 8.32 1.14
                 8.00 1.14 8.00 0.90 7.64 0.90 7.64 1.14 7.32 1.14 7.32 0.90
                 6.24 0.90 6.24 1.14 5.92 1.14 5.92 0.90 4.84 0.90 4.84 1.14
                 4.52 1.14 4.52 0.90 1.28 0.90 1.28 1.58 0.96 1.58 0.96 0.90
                 0.00 0.90 0.00 -0.90 11.52 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 11.52 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  11.16 4.10 10.84 4.10 10.84 1.78 9.66 1.78 9.66 2.65 8.56 2.65
                 8.56 2.33 9.34 2.33 9.34 1.46 10.84 1.46 10.84 1.22 11.16 1.22 ;
        POLYGON  10.37 4.54 0.16 4.54 0.16 1.26 0.50 1.26 0.50 1.58 0.48 1.58
                 0.48 3.10 1.94 3.10 1.94 3.42 0.48 3.42 0.48 4.22 10.05 4.22
                 10.05 2.66 9.98 2.66 9.98 2.34 10.37 2.34 ;
        RECT  8.52 3.58 9.52 3.90 ;
        POLYGON  9.02 1.78 8.24 1.78 8.24 2.34 8.14 2.34 8.14 3.90 7.82 3.90
                 7.82 2.81 7.03 2.81 7.03 2.48 7.82 2.48 7.82 2.02 7.92 2.02
                 7.92 1.46 9.02 1.46 ;
        POLYGON  4.66 3.26 2.58 3.26 2.58 3.90 2.26 3.90 2.26 2.93 3.20 2.93
                 3.20 1.22 3.52 1.22 3.52 2.93 4.66 2.93 ;
        RECT  1.82 1.22 2.84 1.54 ;
    END
END tinvh_16

MACRO tinvh_12
    CLASS CORE ;
    FOREIGN tinvh_12 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.52 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.72 ;
        END
    END a
    PIN en
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.06  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 1.76 2.72 ;
        END
    END en
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.28  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  6.94 1.78 5.60 1.78 5.60 3.58 6.78 3.58 6.78 3.90 3.64 3.90
                 3.64 3.58 5.28 3.58 5.28 1.78 5.22 1.78 5.22 1.46 6.94 1.46 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  11.52 0.90 10.46 0.90 10.46 1.14 10.14 1.14 10.14 0.90
                 9.74 0.90 9.74 1.14 9.42 1.14 9.42 0.90 8.32 0.90 8.32 1.14
                 8.00 1.14 8.00 0.90 7.64 0.90 7.64 1.14 7.32 1.14 7.32 0.90
                 6.24 0.90 6.24 1.14 5.92 1.14 5.92 0.90 4.84 0.90 4.84 1.14
                 4.52 1.14 4.52 0.90 1.28 0.90 1.28 1.58 0.96 1.58 0.96 0.90
                 0.00 0.90 0.00 -0.90 11.52 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 11.52 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  11.16 4.10 10.84 4.10 10.84 1.78 9.66 1.78 9.66 2.65 8.56 2.65
                 8.56 2.33 9.34 2.33 9.34 1.46 10.84 1.46 10.84 1.22 11.16 1.22 ;
        POLYGON  10.37 4.54 0.16 4.54 0.16 1.26 0.50 1.26 0.50 1.58 0.48 1.58
                 0.48 3.10 1.94 3.10 1.94 3.42 0.48 3.42 0.48 4.22 10.05 4.22
                 10.05 2.66 9.98 2.66 9.98 2.34 10.37 2.34 ;
        RECT  8.52 3.58 9.52 3.90 ;
        POLYGON  9.02 1.78 8.24 1.78 8.24 2.34 8.14 2.34 8.14 3.90 7.82 3.90
                 7.82 2.81 7.03 2.81 7.03 2.48 7.82 2.48 7.82 2.02 7.92 2.02
                 7.92 1.46 9.02 1.46 ;
        POLYGON  4.66 3.26 2.58 3.26 2.58 3.90 2.26 3.90 2.26 2.93 3.20 2.93
                 3.20 1.22 3.52 1.22 3.52 2.93 4.66 2.93 ;
        RECT  1.82 1.22 2.84 1.54 ;
    END
END tinvh_12

MACRO tinvh_10
    CLASS CORE ;
    FOREIGN tinvh_10 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.88 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.72 ;
        END
    END a
    PIN en
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.06  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 1.76 2.72 ;
        END
    END en
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.97  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  6.78 3.90 3.64 3.90 3.64 3.58 5.28 3.58 5.28 1.78 4.68 1.78
                 4.68 1.46 6.40 1.46 6.40 1.78 5.60 1.78 5.60 3.58 6.78 3.58 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  10.88 0.90 9.92 0.90 9.92 1.14 9.60 1.14 9.60 0.90 9.20 0.90
                 9.20 1.14 8.88 1.14 8.88 0.90 7.78 0.90 7.78 1.14 7.46 1.14
                 7.46 0.90 7.10 0.90 7.10 1.14 6.78 1.14 6.78 0.90 5.70 0.90
                 5.70 1.14 5.38 1.14 5.38 0.90 4.30 0.90 4.30 1.14 3.98 1.14
                 3.98 0.90 1.28 0.90 1.28 1.58 0.96 1.58 0.96 0.90 0.00 0.90
                 0.00 -0.90 10.88 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 10.88 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  10.62 4.10 10.30 4.10 10.30 1.78 9.12 1.78 9.12 2.65 8.02 2.65
                 8.02 2.33 8.80 2.33 8.80 1.46 10.30 1.46 10.30 1.22 10.62 1.22 ;
        POLYGON  9.83 4.54 0.16 4.54 0.16 1.26 0.50 1.26 0.50 1.58 0.48 1.58
                 0.48 3.10 1.94 3.10 1.94 3.42 0.48 3.42 0.48 4.22 9.51 4.22
                 9.51 2.66 9.44 2.66 9.44 2.34 9.83 2.34 ;
        RECT  7.98 3.58 8.98 3.90 ;
        POLYGON  8.48 1.78 7.70 1.78 7.70 2.34 7.60 2.34 7.60 3.90 7.28 3.90
                 7.28 2.81 6.49 2.81 6.49 2.48 7.28 2.48 7.28 2.02 7.38 2.02
                 7.38 1.46 8.48 1.46 ;
        POLYGON  4.66 3.26 2.58 3.26 2.58 3.90 2.26 3.90 2.26 2.93 3.20 2.93
                 3.20 1.22 3.52 1.22 3.52 2.93 4.66 2.93 ;
        RECT  1.82 1.22 2.84 1.54 ;
    END
END tinvh_10

MACRO tinvh_1
    CLASS CORE ;
    FOREIGN tinvh_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.96 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.45  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.72 ;
        END
    END a
    PIN en
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.02  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 1.76 2.72 ;
        END
    END en
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.39  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  5.19 1.54 5.07 1.54 4.98 1.63 4.98 3.90 4.47 3.90 4.47 3.58
                 4.66 3.58 4.66 2.40 4.64 2.40 4.64 2.08 4.66 2.08 4.66 1.43
                 4.87 1.22 5.19 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.96 0.90 8.08 0.90 8.08 1.14 7.76 1.14 7.76 0.90 7.36 0.90
                 7.36 1.14 7.04 1.14 7.04 0.90 5.87 0.90 5.87 1.14 5.55 1.14
                 5.55 0.90 4.49 0.90 4.49 1.14 4.17 1.14 4.17 0.90 1.28 0.90
                 1.28 1.58 0.96 1.58 0.96 0.90 0.00 0.90 0.00 -0.90 8.96 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 8.96 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  8.78 4.34 8.46 4.34 8.46 1.78 7.21 1.78 7.21 2.65 6.18 2.65
                 6.18 2.33 6.89 2.33 6.89 1.46 8.46 1.46 8.46 1.22 8.78 1.22 ;
        POLYGON  7.99 4.54 0.16 4.54 0.16 1.26 0.50 1.26 0.50 1.58 0.48 1.58
                 0.48 3.10 1.94 3.10 1.94 3.42 0.48 3.42 0.48 4.22 7.67 4.22
                 7.67 2.66 7.56 2.66 7.56 2.34 7.99 2.34 ;
        RECT  6.14 3.58 7.14 3.90 ;
        POLYGON  6.57 1.78 5.86 1.78 5.86 2.34 5.76 2.34 5.76 3.90 5.44 3.90
                 5.44 2.34 5.30 2.34 5.30 2.02 5.54 2.02 5.54 1.46 6.57 1.46 ;
        POLYGON  4.34 2.96 2.58 2.96 2.58 3.90 2.26 3.90 2.26 2.64 3.20 2.64
                 3.20 1.22 3.52 1.22 3.52 2.64 4.34 2.64 ;
        RECT  1.82 1.22 2.84 1.54 ;
    END
END tinvh_1

MACRO tinvh_0
    CLASS CORE ;
    FOREIGN tinvh_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.96 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.45  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.72 ;
        END
    END a
    PIN en
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.02  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 1.76 2.72 ;
        END
    END en
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.35  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  5.19 1.54 5.07 1.54 4.98 1.63 4.98 3.90 4.47 3.90 4.47 3.58
                 4.66 3.58 4.66 2.40 4.64 2.40 4.64 2.08 4.66 2.08 4.66 1.43
                 4.87 1.22 5.19 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.96 0.90 8.08 0.90 8.08 1.14 7.76 1.14 7.76 0.90 7.36 0.90
                 7.36 1.14 7.04 1.14 7.04 0.90 5.87 0.90 5.87 1.14 5.55 1.14
                 5.55 0.90 4.49 0.90 4.49 1.14 4.17 1.14 4.17 0.90 1.28 0.90
                 1.28 1.58 0.96 1.58 0.96 0.90 0.00 0.90 0.00 -0.90 8.96 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 8.96 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  8.78 4.34 8.46 4.34 8.46 1.78 7.21 1.78 7.21 2.65 6.18 2.65
                 6.18 2.33 6.89 2.33 6.89 1.46 8.46 1.46 8.46 1.22 8.78 1.22 ;
        POLYGON  7.99 4.54 0.16 4.54 0.16 1.26 0.50 1.26 0.50 1.58 0.48 1.58
                 0.48 3.10 1.94 3.10 1.94 3.42 0.48 3.42 0.48 4.22 7.67 4.22
                 7.67 2.66 7.56 2.66 7.56 2.34 7.99 2.34 ;
        RECT  6.14 3.58 7.14 3.90 ;
        POLYGON  6.57 1.78 5.86 1.78 5.86 2.34 5.76 2.34 5.76 3.90 5.44 3.90
                 5.44 2.34 5.30 2.34 5.30 2.02 5.54 2.02 5.54 1.46 6.57 1.46 ;
        POLYGON  4.34 2.96 2.58 2.96 2.58 3.90 2.26 3.90 2.26 2.64 3.20 2.64
                 3.20 1.22 3.52 1.22 3.52 2.64 4.34 2.64 ;
        RECT  1.82 1.22 2.84 1.54 ;
    END
END tinvh_0

MACRO tielo
    CLASS CORE TIELOW ;
    FOREIGN tielo 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 1.92 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 1.38 1.76 1.76 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  1.92 0.90 0.74 0.90 0.74 1.32 0.42 1.32 0.42 0.90 0.00 0.90
                 0.00 -0.90 1.92 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  1.92 6.66 0.00 6.66 0.00 4.86 0.42 4.86 0.42 3.40 0.74 3.40
                 0.74 4.86 1.92 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  1.44 4.34 1.12 4.34 1.12 2.56 0.80 2.56 0.80 2.24 1.44 2.24 ;
    END
END tielo

MACRO tiehi
    CLASS CORE TIEHIGH ;
    FOREIGN tiehi 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 1.92 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.70  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.76 3.68 1.44 3.68 1.44 4.34 1.12 4.34 1.12 3.36 1.76 3.36 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  1.92 0.90 0.74 0.90 0.74 1.32 0.42 1.32 0.42 0.90 0.00 0.90
                 0.00 -0.90 1.92 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  1.92 6.66 0.00 6.66 0.00 4.86 0.42 4.86 0.42 3.40 0.74 3.40
                 0.74 4.86 1.92 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  1.44 1.96 1.12 1.96 1.12 2.56 0.80 2.56 0.80 1.64 1.12 1.64
                 1.12 1.38 1.44 1.38 ;
    END
END tiehi

MACRO tbufh_8
    CLASS CORE ;
    FOREIGN tbufh_8 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.60 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.23  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.57 4.54 0.80 4.54 0.80 3.10 1.24 3.10 1.24 3.42 1.12 3.42
                 1.12 4.22 8.25 4.22 8.25 2.66 8.18 2.66 8.18 2.34 8.57 2.34 ;
        END
    END a
    PIN en
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.06  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.74 2.08 1.12 2.72 ;
        END
    END en
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.74  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  5.14 1.54 5.02 1.54 4.96 1.60 4.96 3.90 2.94 3.90 2.94 3.58
                 4.64 3.58 4.64 1.40 4.82 1.22 5.14 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  9.60 0.90 8.66 0.90 8.66 1.14 8.34 1.14 8.34 0.90 7.94 0.90
                 7.94 1.14 7.62 1.14 7.62 0.90 6.52 0.90 6.52 1.14 6.20 1.14
                 6.20 0.90 5.84 0.90 5.84 1.14 5.52 1.14 5.52 0.90 4.44 0.90
                 4.44 1.14 4.12 1.14 4.12 0.90 0.74 0.90 0.74 1.58 0.42 1.58
                 0.42 0.90 0.00 0.90 0.00 -0.90 9.60 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 9.60 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  9.36 4.10 9.04 4.10 9.04 1.78 7.86 1.78 7.86 2.65 6.76 2.65
                 6.76 2.33 7.54 2.33 7.54 1.46 9.04 1.46 9.04 1.22 9.36 1.22 ;
        RECT  6.72 3.58 7.72 3.90 ;
        POLYGON  7.22 1.78 6.44 1.78 6.44 2.34 6.34 2.34 6.34 3.90 6.02 3.90
                 6.02 2.98 5.39 2.98 5.39 2.66 6.02 2.66 6.02 2.02 6.12 2.02
                 6.12 1.46 7.22 1.46 ;
        POLYGON  3.76 2.89 1.88 2.89 1.88 3.90 1.56 3.90 1.56 2.57 2.50 2.57
                 2.50 1.22 2.82 1.22 2.82 2.57 3.76 2.57 ;
        RECT  1.12 1.22 2.14 1.54 ;
    END
END tbufh_8

MACRO tbufh_64
    CLASS CORE ;
    FOREIGN tbufh_64 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 31.36 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 4.94  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  23.31 2.60 22.68 2.60 22.68 3.67 21.61 3.67 21.61 4.53
                 21.54 4.53 21.54 4.54 0.16 4.54 0.16 2.90 2.50 2.90 2.50 3.22
                 0.48 3.22 0.48 4.22 21.29 4.22 21.29 3.35 22.36 3.35
                 22.36 2.28 23.31 2.28 ;
        END
    END a
    PIN en
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  7.79 1.80 8.16 2.62 ;
        END
    END en
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 16.39  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.88 3.90 17.65 3.90 17.65 1.78 15.30 1.78 15.30 3.58
                 17.65 3.58 17.65 3.90 14.98 3.90 14.98 1.78 12.64 1.78
                 12.64 3.58 14.98 3.58 14.98 3.90 12.32 3.90 12.32 1.78
                 9.70 1.78 9.70 3.58 12.32 3.58 12.32 3.90 7.91 3.90 7.91 3.58
                 9.38 3.58 9.38 1.46 19.50 1.46 19.50 1.78 17.97 1.78
                 17.97 3.58 20.88 3.58 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  31.36 0.90 29.91 0.90 29.91 1.16 29.59 1.16 29.59 0.90
                 27.49 0.90 27.49 1.16 27.17 1.16 27.17 0.90 26.09 0.90
                 26.09 1.16 25.77 1.16 25.77 0.90 24.69 0.90 24.69 1.16
                 24.37 1.16 24.37 0.90 23.29 0.90 23.29 1.16 22.97 1.16
                 22.97 0.90 20.20 0.90 20.20 1.14 19.88 1.14 19.88 0.90
                 18.80 0.90 18.80 1.14 18.48 1.14 18.48 0.90 17.40 0.90
                 17.40 1.14 17.08 1.14 17.08 0.90 16.00 0.90 16.00 1.14
                 15.68 1.14 15.68 0.90 14.60 0.90 14.60 1.14 14.28 1.14
                 14.28 0.90 13.20 0.90 13.20 1.14 12.88 1.14 12.88 0.90
                 11.80 0.90 11.80 1.14 11.48 1.14 11.48 0.90 10.40 0.90
                 10.40 1.14 10.08 1.14 10.08 0.90 9.00 0.90 9.00 1.14 8.68 1.14
                 8.68 0.90 0.00 0.90 0.00 -0.90 31.36 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 31.36 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  30.61 1.80 29.21 1.80 29.21 3.43 30.61 3.43 30.61 4.54
                 30.29 4.54 30.29 3.75 29.21 3.75 29.21 4.54 28.89 4.54
                 28.89 2.62 26.87 2.62 26.87 2.30 28.89 2.30 28.89 1.48
                 30.61 1.48 ;
        POLYGON  28.53 3.85 28.21 3.85 28.21 3.26 27.13 3.26 27.13 3.85
                 26.81 3.85 26.81 3.26 25.73 3.26 25.73 3.85 25.41 3.85
                 25.41 1.92 21.79 1.92 21.79 2.81 18.80 2.81 18.80 2.48
                 21.47 2.48 21.47 1.60 28.19 1.60 28.19 1.92 25.73 1.92
                 25.73 2.94 28.53 2.94 ;
        RECT  21.93 4.17 27.87 4.49 ;
        POLYGON  8.86 3.26 6.72 3.26 6.72 3.90 0.80 3.90 0.80 3.58 6.40 3.58
                 6.40 2.34 4.28 2.34 4.28 2.02 7.08 2.02 7.08 1.34 7.40 1.34
                 7.40 2.34 6.72 2.34 6.72 2.94 8.86 2.94 ;
        RECT  0.80 1.32 6.70 1.64 ;
    END
END tbufh_64

MACRO tbufh_6
    CLASS CORE ;
    FOREIGN tbufh_6 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.60 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.23  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.57 4.54 0.80 4.54 0.80 3.10 1.24 3.10 1.24 3.42 1.12 3.42
                 1.12 4.22 8.25 4.22 8.25 2.66 8.18 2.66 8.18 2.34 8.57 2.34 ;
        END
    END a
    PIN en
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.06  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.74 2.08 1.12 2.72 ;
        END
    END en
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.62  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  5.14 1.54 5.02 1.54 4.96 1.60 4.96 3.90 2.94 3.90 2.94 3.58
                 4.64 3.58 4.64 1.40 4.82 1.22 5.14 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  9.60 0.90 8.66 0.90 8.66 1.14 8.34 1.14 8.34 0.90 7.94 0.90
                 7.94 1.14 7.62 1.14 7.62 0.90 6.52 0.90 6.52 1.14 6.20 1.14
                 6.20 0.90 5.84 0.90 5.84 1.14 5.52 1.14 5.52 0.90 4.44 0.90
                 4.44 1.14 4.12 1.14 4.12 0.90 0.74 0.90 0.74 1.58 0.42 1.58
                 0.42 0.90 0.00 0.90 0.00 -0.90 9.60 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 9.60 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  9.36 4.10 9.04 4.10 9.04 1.78 7.86 1.78 7.86 2.65 6.76 2.65
                 6.76 2.33 7.54 2.33 7.54 1.46 9.04 1.46 9.04 1.22 9.36 1.22 ;
        RECT  6.72 3.58 7.72 3.90 ;
        POLYGON  7.22 1.78 6.44 1.78 6.44 2.34 6.34 2.34 6.34 3.90 6.02 3.90
                 6.02 2.98 5.28 2.98 5.28 2.66 6.02 2.66 6.02 2.02 6.12 2.02
                 6.12 1.46 7.22 1.46 ;
        POLYGON  3.76 2.89 1.88 2.89 1.88 3.90 1.56 3.90 1.56 2.57 2.50 2.57
                 2.50 1.22 2.82 1.22 2.82 2.57 3.76 2.57 ;
        RECT  1.12 1.22 2.14 1.54 ;
    END
END tbufh_6

MACRO tbufh_48
    CLASS CORE ;
    FOREIGN tbufh_48 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 30.72 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 4.94  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  23.31 2.60 22.68 2.60 22.68 3.67 21.61 3.67 21.61 4.53
                 21.54 4.53 21.54 4.54 0.16 4.54 0.16 2.90 2.50 2.90 2.50 3.22
                 0.48 3.22 0.48 4.22 21.29 4.22 21.29 3.35 22.36 3.35
                 22.36 2.28 23.31 2.28 ;
        END
    END a
    PIN en
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.97  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  7.79 1.86 8.16 2.62 ;
        END
    END en
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 15.82  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.88 3.90 17.65 3.90 17.65 1.78 15.30 1.78 15.30 3.58
                 17.65 3.58 17.65 3.90 14.98 3.90 14.98 1.78 12.00 1.78
                 12.00 3.58 14.98 3.58 14.98 3.90 11.68 3.90 11.68 1.78
                 9.70 1.78 9.70 3.58 11.68 3.58 11.68 3.90 7.91 3.90 7.91 3.58
                 9.38 3.58 9.38 1.46 19.50 1.46 19.50 1.78 17.97 1.78
                 17.97 3.58 20.88 3.58 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  30.72 0.90 29.21 0.90 29.21 1.16 28.89 1.16 28.89 0.90
                 27.49 0.90 27.49 1.16 27.17 1.16 27.17 0.90 26.09 0.90
                 26.09 1.16 25.77 1.16 25.77 0.90 24.69 0.90 24.69 1.16
                 24.37 1.16 24.37 0.90 23.29 0.90 23.29 1.16 22.97 1.16
                 22.97 0.90 20.20 0.90 20.20 1.14 19.88 1.14 19.88 0.90
                 18.80 0.90 18.80 1.14 18.48 1.14 18.48 0.90 17.40 0.90
                 17.40 1.14 17.08 1.14 17.08 0.90 16.00 0.90 16.00 1.14
                 15.68 1.14 15.68 0.90 14.60 0.90 14.60 1.14 14.28 1.14
                 14.28 0.90 13.20 0.90 13.20 1.14 12.88 1.14 12.88 0.90
                 11.80 0.90 11.80 1.14 11.48 1.14 11.48 0.90 10.40 0.90
                 10.40 1.14 10.08 1.14 10.08 0.90 9.00 0.90 9.00 1.14 8.68 1.14
                 8.68 0.90 0.00 0.90 0.00 -0.90 30.72 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 30.72 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  29.91 4.54 29.59 4.54 29.59 2.62 26.87 2.62 26.87 2.30
                 29.59 2.30 29.59 1.48 29.91 1.48 ;
        POLYGON  28.53 3.85 28.21 3.85 28.21 3.26 27.13 3.26 27.13 3.85
                 26.81 3.85 26.81 3.26 25.73 3.26 25.73 3.85 25.41 3.85
                 25.41 1.92 21.79 1.92 21.79 2.81 18.80 2.81 18.80 2.48
                 21.47 2.48 21.47 1.60 28.19 1.60 28.19 1.92 25.73 1.92
                 25.73 2.94 28.53 2.94 ;
        RECT  21.93 4.17 27.87 4.49 ;
        POLYGON  8.86 3.26 6.72 3.26 6.72 3.90 0.80 3.90 0.80 3.58 6.40 3.58
                 6.40 2.34 4.28 2.34 4.28 2.02 7.08 2.02 7.08 1.34 7.40 1.34
                 7.40 2.34 6.72 2.34 6.72 2.94 8.86 2.94 ;
        RECT  0.80 1.32 6.70 1.64 ;
    END
END tbufh_48

MACRO tbufh_4
    CLASS CORE ;
    FOREIGN tbufh_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.32 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.23  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.29 4.54 0.80 4.54 0.80 3.10 1.24 3.10 1.24 3.42 1.12 3.42
                 1.12 4.22 6.97 4.22 6.97 2.66 6.86 2.66 6.86 2.34 7.29 2.34 ;
        END
    END a
    PIN en
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.06  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.74 2.08 1.12 2.72 ;
        END
    END en
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.64  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.49 1.54 4.37 1.54 4.28 1.63 4.28 2.72 4.32 2.72 4.32 3.90
                 3.69 3.90 3.69 3.58 4.00 3.58 4.00 3.04 3.96 3.04 3.96 1.43
                 4.17 1.22 4.49 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 0.90 7.38 0.90 7.38 1.14 7.06 1.14 7.06 0.90 6.66 0.90
                 6.66 1.14 6.34 1.14 6.34 0.90 5.17 0.90 5.17 1.14 4.85 1.14
                 4.85 0.90 3.79 0.90 3.79 1.14 3.47 1.14 3.47 0.90 0.74 0.90
                 0.74 1.58 0.42 1.58 0.42 0.90 0.00 0.90 0.00 -0.90 8.32 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 8.32 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  8.08 4.10 7.76 4.10 7.76 1.78 6.51 1.78 6.51 2.65 5.48 2.65
                 5.48 2.33 6.19 2.33 6.19 1.46 7.76 1.46 7.76 1.22 8.08 1.22 ;
        RECT  5.44 3.58 6.44 3.90 ;
        POLYGON  5.87 1.78 5.16 1.78 5.16 2.34 5.06 2.34 5.06 3.90 4.74 3.90
                 4.74 2.34 4.60 2.34 4.60 2.02 4.84 2.02 4.84 1.46 5.87 1.46 ;
        POLYGON  3.64 2.96 1.88 2.96 1.88 3.90 1.56 3.90 1.56 2.64 2.50 2.64
                 2.50 1.22 2.82 1.22 2.82 2.64 3.64 2.64 ;
        RECT  1.12 1.22 2.14 1.54 ;
    END
END tbufh_4

MACRO tbufh_32
    CLASS CORE ;
    FOREIGN tbufh_32 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 17.28 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.47  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.29 4.54 0.16 4.54 0.16 2.94 1.26 2.94 1.26 3.26 0.48 3.26
                 0.48 4.22 15.97 4.22 15.97 3.26 13.94 3.26 13.94 2.94
                 16.29 2.94 ;
        END
    END a
    PIN en
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.83  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.86 1.14 2.48 ;
        END
    END en
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 8.89  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  11.74 3.90 9.15 3.90 9.15 1.78 6.88 1.78 6.88 3.58 9.15 3.58
                 9.15 3.90 4.42 3.90 4.42 3.58 6.56 3.58 6.56 1.78 6.00 1.78
                 6.00 1.46 10.52 1.46 10.52 1.78 9.47 1.78 9.47 3.58 11.74 3.58 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  17.28 0.90 14.84 0.90 14.84 1.14 14.52 1.14 14.52 0.90
                 13.44 0.90 13.44 1.14 13.12 1.14 13.12 0.90 11.22 0.90
                 11.22 1.14 10.90 1.14 10.90 0.90 9.82 0.90 9.82 1.14 9.50 1.14
                 9.50 0.90 8.42 0.90 8.42 1.14 8.10 1.14 8.10 0.90 7.02 0.90
                 7.02 1.14 6.70 1.14 6.70 0.90 5.62 0.90 5.62 1.14 5.30 1.14
                 5.30 0.90 0.74 0.90 0.74 1.54 0.42 1.54 0.42 0.90 0.00 0.90
                 0.00 -0.90 17.28 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 17.28 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  17.08 4.10 16.76 4.10 16.76 2.62 13.48 2.62 13.48 2.30
                 16.76 2.30 16.76 1.22 17.08 1.22 ;
        POLYGON  15.54 1.78 13.14 1.78 13.14 3.26 12.80 3.26 12.80 2.80
                 9.92 2.80 9.92 2.48 12.80 2.48 12.80 1.78 12.42 1.78
                 12.42 1.46 15.54 1.46 ;
        RECT  12.10 3.58 15.40 3.90 ;
        POLYGON  6.14 3.26 4.06 3.26 4.06 3.90 3.74 3.90 3.74 3.26 2.66 3.26
                 2.66 3.90 0.94 3.90 0.94 3.58 2.34 3.58 2.34 2.94 3.28 2.94
                 3.28 1.86 3.60 1.86 3.60 2.94 6.14 2.94 ;
        RECT  1.20 1.22 4.30 1.54 ;
    END
END tbufh_32

MACRO tbufh_3
    CLASS CORE ;
    FOREIGN tbufh_3 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.32 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.23  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.29 4.54 0.80 4.54 0.80 3.07 1.24 3.07 1.24 3.71 1.12 3.71
                 1.12 4.22 6.97 4.22 6.97 2.66 6.86 2.66 6.86 2.34 7.29 2.34 ;
        END
    END a
    PIN en
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.02  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.74 2.08 1.12 2.72 ;
        END
    END en
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.49 1.54 4.37 1.54 4.28 1.63 4.28 2.72 4.32 2.72 4.32 3.90
                 3.69 3.90 3.69 3.58 4.00 3.58 4.00 3.04 3.96 3.04 3.96 1.43
                 4.17 1.22 4.49 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 0.90 7.38 0.90 7.38 1.14 7.06 1.14 7.06 0.90 6.66 0.90
                 6.66 1.14 6.34 1.14 6.34 0.90 5.17 0.90 5.17 1.14 4.85 1.14
                 4.85 0.90 3.79 0.90 3.79 1.14 3.47 1.14 3.47 0.90 0.74 0.90
                 0.74 1.58 0.42 1.58 0.42 0.90 0.00 0.90 0.00 -0.90 8.32 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 8.32 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  8.08 4.34 7.76 4.34 7.76 1.78 6.51 1.78 6.51 2.65 5.48 2.65
                 5.48 2.33 6.19 2.33 6.19 1.46 7.76 1.46 7.76 1.22 8.08 1.22 ;
        RECT  5.44 3.58 6.44 3.90 ;
        POLYGON  5.87 1.78 5.16 1.78 5.16 2.34 5.06 2.34 5.06 3.90 4.74 3.90
                 4.74 2.34 4.60 2.34 4.60 2.02 4.84 2.02 4.84 1.46 5.87 1.46 ;
        POLYGON  3.64 2.96 1.88 2.96 1.88 3.90 1.56 3.90 1.56 2.64 2.50 2.64
                 2.50 1.22 2.82 1.22 2.82 2.64 3.64 2.64 ;
        RECT  1.12 1.22 2.14 1.54 ;
    END
END tbufh_3

MACRO tbufh_24
    CLASS CORE ;
    FOREIGN tbufh_24 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 17.28 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.47  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.21 4.54 0.16 4.54 0.16 2.94 1.18 2.94 1.18 3.26 0.48 3.26
                 0.48 4.22 15.89 4.22 15.89 3.26 13.86 3.26 13.86 2.94
                 16.21 2.94 ;
        END
    END a
    PIN en
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.83  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.74 1.86 1.12 2.48 ;
        END
    END en
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 8.56  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  11.66 3.90 9.07 3.90 9.07 1.78 6.88 1.78 6.88 3.58 9.07 3.58
                 9.07 3.90 4.34 3.90 4.34 3.58 6.56 3.58 6.56 1.78 5.92 1.78
                 5.92 1.46 10.44 1.46 10.44 1.78 9.39 1.78 9.39 3.58 11.66 3.58 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  17.28 0.90 14.76 0.90 14.76 1.14 14.44 1.14 14.44 0.90
                 13.36 0.90 13.36 1.14 13.04 1.14 13.04 0.90 11.14 0.90
                 11.14 1.14 10.82 1.14 10.82 0.90 9.74 0.90 9.74 1.14 9.42 1.14
                 9.42 0.90 8.34 0.90 8.34 1.14 8.02 1.14 8.02 0.90 6.94 0.90
                 6.94 1.14 6.62 1.14 6.62 0.90 5.54 0.90 5.54 1.14 5.22 1.14
                 5.22 0.90 0.74 0.90 0.74 1.54 0.42 1.54 0.42 0.90 0.00 0.90
                 0.00 -0.90 17.28 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 17.28 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  17.00 4.10 16.68 4.10 16.68 2.62 13.40 2.62 13.40 2.30
                 16.68 2.30 16.68 1.22 17.00 1.22 ;
        POLYGON  15.46 1.78 13.06 1.78 13.06 3.26 12.72 3.26 12.72 2.80
                 9.84 2.80 9.84 2.48 12.72 2.48 12.72 1.78 12.34 1.78
                 12.34 1.46 15.46 1.46 ;
        RECT  12.02 3.58 15.32 3.90 ;
        POLYGON  6.06 3.26 3.98 3.26 3.98 3.90 3.66 3.90 3.66 3.26 2.58 3.26
                 2.58 3.90 0.86 3.90 0.86 3.58 2.26 3.58 2.26 2.94 3.20 2.94
                 3.20 1.86 3.52 1.86 3.52 2.94 6.06 2.94 ;
        RECT  1.12 1.22 4.22 1.54 ;
    END
END tbufh_24

MACRO tbufh_20
    CLASS CORE ;
    FOREIGN tbufh_20 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.00 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.47  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  15.01 4.54 0.16 4.54 0.16 2.94 1.26 2.94 1.26 3.26 0.48 3.26
                 0.48 4.22 14.69 4.22 14.69 3.26 12.66 3.26 12.66 2.94
                 15.01 2.94 ;
        END
    END a
    PIN en
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.86 1.14 2.48 ;
        END
    END en
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 7.22  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.34 3.90 8.28 3.90 8.28 1.78 6.88 1.78 6.88 3.58 8.28 3.58
                 8.28 3.90 4.42 3.90 4.42 3.58 6.56 3.58 6.56 1.78 5.46 1.78
                 5.46 1.46 9.98 1.46 9.98 1.78 8.60 1.78 8.60 3.58 10.34 3.58 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 0.90 13.56 0.90 13.56 1.14 13.24 1.14 13.24 0.90
                 12.16 0.90 12.16 1.14 11.84 1.14 11.84 0.90 10.68 0.90
                 10.68 1.14 10.36 1.14 10.36 0.90 9.28 0.90 9.28 1.14 8.96 1.14
                 8.96 0.90 7.88 0.90 7.88 1.14 7.56 1.14 7.56 0.90 6.48 0.90
                 6.48 1.14 6.16 1.14 6.16 0.90 5.08 0.90 5.08 1.14 4.76 1.14
                 4.76 0.90 0.00 0.90 0.00 -0.90 16.00 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 16.00 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  15.80 4.39 15.48 4.39 15.48 2.62 12.20 2.62 12.20 2.30
                 15.48 2.30 15.48 1.22 15.80 1.22 ;
        POLYGON  14.26 1.78 11.86 1.78 11.86 3.26 11.52 3.26 11.52 2.80
                 9.38 2.80 9.38 2.48 11.52 2.48 11.52 1.78 11.14 1.78
                 11.14 1.46 14.26 1.46 ;
        RECT  10.82 3.58 14.12 3.90 ;
        POLYGON  6.15 3.26 4.06 3.26 4.06 3.90 3.74 3.90 3.74 3.26 2.66 3.26
                 2.66 3.90 0.94 3.90 0.94 3.58 2.34 3.58 2.34 2.94 3.28 2.94
                 3.28 1.86 3.60 1.86 3.60 2.94 6.15 2.94 ;
        RECT  1.20 1.22 4.30 1.54 ;
    END
END tbufh_20

MACRO tbufh_2
    CLASS CORE ;
    FOREIGN tbufh_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.32 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.23  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.29 4.54 0.80 4.54 0.80 3.10 1.24 3.10 1.24 4.22 6.97 4.22
                 6.97 2.66 6.86 2.66 6.86 2.34 7.29 2.34 ;
        END
    END a
    PIN en
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.02  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.12 2.40 1.06 2.40 1.06 2.72 0.74 2.72 0.74 2.08 1.12 2.08 ;
        END
    END en
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.38  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.49 1.54 4.37 1.54 4.28 1.63 4.28 2.72 4.32 2.72 4.32 3.90
                 3.69 3.90 3.69 3.58 4.00 3.58 4.00 3.04 3.96 3.04 3.96 2.40
                 3.94 2.40 3.94 2.08 3.96 2.08 3.96 1.43 4.17 1.22 4.49 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 0.90 7.38 0.90 7.38 1.14 7.06 1.14 7.06 0.90 6.66 0.90
                 6.66 1.14 6.34 1.14 6.34 0.90 5.17 0.90 5.17 1.14 4.85 1.14
                 4.85 0.90 3.79 0.90 3.79 1.14 3.47 1.14 3.47 0.90 0.74 0.90
                 0.74 1.58 0.42 1.58 0.42 0.90 0.00 0.90 0.00 -0.90 8.32 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 8.32 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  8.08 4.34 7.76 4.34 7.76 1.78 6.51 1.78 6.51 2.65 5.48 2.65
                 5.48 2.33 6.19 2.33 6.19 1.46 7.76 1.46 7.76 1.22 8.08 1.22 ;
        RECT  5.44 3.58 6.44 3.90 ;
        POLYGON  5.87 1.78 5.16 1.78 5.16 2.34 5.06 2.34 5.06 3.90 4.74 3.90
                 4.74 2.34 4.60 2.34 4.60 2.02 4.84 2.02 4.84 1.46 5.87 1.46 ;
        POLYGON  3.64 2.96 1.88 2.96 1.88 3.90 1.56 3.90 1.56 2.64 2.50 2.64
                 2.50 1.22 2.82 1.22 2.82 2.64 3.64 2.64 ;
        RECT  1.12 1.22 2.14 1.54 ;
    END
END tbufh_2

MACRO tbufh_16
    CLASS CORE ;
    FOREIGN tbufh_16 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.88 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.23  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.39 3.61 6.36 3.61 6.36 4.54 0.46 4.54 0.46 2.53 1.14 2.53
                 1.14 3.04 0.80 3.04 0.80 4.22 6.04 4.22 6.04 3.29 7.07 3.29
                 7.07 2.28 7.39 2.28 ;
        END
    END a
    PIN en
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.06  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 1.96 3.18 2.62 ;
        END
    END en
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.44  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  5.80 2.12 4.32 2.12 4.32 3.58 5.62 3.58 5.62 3.90 2.50 3.90
                 2.50 3.58 4.00 3.58 4.00 1.80 5.80 1.80 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  10.88 0.90 9.76 0.90 9.76 1.58 9.44 1.58 9.44 0.90 8.04 0.90
                 8.04 1.16 7.72 1.16 7.72 0.90 6.50 0.90 6.50 1.16 6.18 1.16
                 6.18 0.90 5.10 0.90 5.10 1.16 4.78 1.16 4.78 0.92 3.70 0.92
                 3.70 1.16 3.38 1.16 3.38 0.90 0.00 0.90 0.00 -0.90 10.88 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 10.88 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  10.46 4.42 10.14 4.42 10.14 2.62 8.35 2.62 8.35 2.30
                 10.14 2.30 10.14 1.48 10.46 1.48 ;
        POLYGON  9.08 3.85 8.76 3.85 8.76 3.26 7.71 3.26 7.71 1.92 6.72 1.92
                 6.72 2.82 4.77 2.82 4.77 2.50 6.40 2.50 6.40 1.60 8.74 1.60
                 8.74 1.92 8.03 1.92 8.03 2.94 9.08 2.94 ;
        RECT  6.68 4.17 8.41 4.49 ;
        POLYGON  3.44 3.26 1.90 3.26 1.90 3.90 1.12 3.90 1.12 3.58 1.57 3.58
                 1.57 2.34 1.56 2.34 1.56 2.02 1.90 2.02 1.90 2.94 3.44 2.94 ;
        RECT  0.18 1.32 2.61 1.64 ;
    END
END tbufh_16

MACRO tbufh_12
    CLASS CORE ;
    FOREIGN tbufh_12 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.88 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.28  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  6.24 1.78 4.96 1.78 4.96 3.58 6.08 3.58 6.08 3.90 2.94 3.90
                 2.94 3.58 4.64 3.58 4.64 1.78 4.52 1.78 4.52 1.46 6.24 1.46 ;
        END
    END x
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.23  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.67 4.54 0.80 4.54 0.80 3.10 1.24 3.10 1.24 3.42 1.12 3.42
                 1.12 4.22 9.35 4.22 9.35 2.66 9.28 2.66 9.28 2.34 9.67 2.34 ;
        END
    END a
    PIN en
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.06  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.74 2.08 1.12 2.72 ;
        END
    END en
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  10.88 0.90 9.76 0.90 9.76 1.14 9.44 1.14 9.44 0.90 9.04 0.90
                 9.04 1.14 8.72 1.14 8.72 0.90 7.62 0.90 7.62 1.14 7.30 1.14
                 7.30 0.90 6.94 0.90 6.94 1.14 6.62 1.14 6.62 0.90 5.54 0.90
                 5.54 1.14 5.22 1.14 5.22 0.90 4.14 0.90 4.14 1.14 3.82 1.14
                 3.82 0.90 0.74 0.90 0.74 1.58 0.42 1.58 0.42 0.90 0.00 0.90
                 0.00 -0.90 10.88 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 10.88 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  10.46 4.10 10.14 4.10 10.14 1.78 8.96 1.78 8.96 2.65 7.86 2.65
                 7.86 2.33 8.64 2.33 8.64 1.46 10.14 1.46 10.14 1.22 10.46 1.22 ;
        RECT  7.82 3.58 8.82 3.90 ;
        POLYGON  8.32 1.78 7.54 1.78 7.54 2.34 7.44 2.34 7.44 3.90 7.12 3.90
                 7.12 2.81 6.33 2.81 6.33 2.48 7.12 2.48 7.12 2.02 7.22 2.02
                 7.22 1.46 8.32 1.46 ;
        POLYGON  3.96 3.26 1.88 3.26 1.88 3.90 1.56 3.90 1.56 2.93 2.50 2.93
                 2.50 1.22 2.82 1.22 2.82 2.93 3.96 2.93 ;
        RECT  1.12 1.22 2.14 1.54 ;
    END
END tbufh_12

MACRO tbufh_10
    CLASS CORE ;
    FOREIGN tbufh_10 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.24 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.23  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.13 4.54 0.80 4.54 0.80 3.10 1.24 3.10 1.24 3.42 1.12 3.42
                 1.12 4.22 8.81 4.22 8.81 2.66 8.74 2.66 8.74 2.34 9.13 2.34 ;
        END
    END a
    PIN en
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.06  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.74 2.08 1.12 2.72 ;
        END
    END en
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.97  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  6.08 3.90 2.94 3.90 2.94 3.58 4.64 3.58 4.64 1.78 3.98 1.78
                 3.98 1.46 5.70 1.46 5.70 1.78 4.96 1.78 4.96 3.58 6.08 3.58 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  10.24 0.90 9.22 0.90 9.22 1.14 8.90 1.14 8.90 0.90 8.50 0.90
                 8.50 1.14 8.18 1.14 8.18 0.90 7.08 0.90 7.08 1.14 6.76 1.14
                 6.76 0.90 6.40 0.90 6.40 1.14 6.08 1.14 6.08 0.90 5.00 0.90
                 5.00 1.14 4.68 1.14 4.68 0.90 3.60 0.90 3.60 1.14 3.28 1.14
                 3.28 0.90 0.74 0.90 0.74 1.58 0.42 1.58 0.42 0.90 0.00 0.90
                 0.00 -0.90 10.24 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 10.24 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  9.92 4.10 9.60 4.10 9.60 1.78 8.42 1.78 8.42 2.65 7.32 2.65
                 7.32 2.33 8.10 2.33 8.10 1.46 9.60 1.46 9.60 1.22 9.92 1.22 ;
        RECT  7.28 3.58 8.28 3.90 ;
        POLYGON  7.78 1.78 7.00 1.78 7.00 2.34 6.90 2.34 6.90 3.90 6.58 3.90
                 6.58 2.81 5.79 2.81 5.79 2.48 6.58 2.48 6.58 2.02 6.68 2.02
                 6.68 1.46 7.78 1.46 ;
        POLYGON  3.96 3.26 1.88 3.26 1.88 3.90 1.56 3.90 1.56 2.93 2.50 2.93
                 2.50 1.22 2.82 1.22 2.82 2.93 3.96 2.93 ;
        RECT  1.12 1.22 2.14 1.54 ;
    END
END tbufh_10

MACRO tbufh_1
    CLASS CORE ;
    FOREIGN tbufh_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.32 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.23  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.29 4.54 0.80 4.54 0.80 3.10 1.24 3.10 1.24 4.22 6.97 4.22
                 6.97 2.66 6.86 2.66 6.86 2.34 7.29 2.34 ;
        END
    END a
    PIN en
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.02  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.12 2.40 1.06 2.40 1.06 2.72 0.74 2.72 0.74 2.08 1.12 2.08 ;
        END
    END en
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.49 1.54 4.37 1.54 4.28 1.63 4.28 2.72 4.32 2.72 4.32 3.90
                 3.69 3.90 3.69 3.58 4.00 3.58 4.00 3.04 3.96 3.04 3.96 2.40
                 3.94 2.40 3.94 2.08 3.96 2.08 3.96 1.43 4.17 1.22 4.49 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 0.90 7.38 0.90 7.38 1.14 7.06 1.14 7.06 0.90 6.66 0.90
                 6.66 1.14 6.34 1.14 6.34 0.90 5.17 0.90 5.17 1.14 4.85 1.14
                 4.85 0.90 3.79 0.90 3.79 1.14 3.47 1.14 3.47 0.90 0.74 0.90
                 0.74 1.58 0.42 1.58 0.42 0.90 0.00 0.90 0.00 -0.90 8.32 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 8.32 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  8.08 4.34 7.76 4.34 7.76 1.78 6.51 1.78 6.51 2.65 5.48 2.65
                 5.48 2.33 6.19 2.33 6.19 1.46 7.76 1.46 7.76 1.22 8.08 1.22 ;
        RECT  5.44 3.58 6.44 3.90 ;
        POLYGON  5.87 1.78 5.16 1.78 5.16 2.34 5.06 2.34 5.06 3.90 4.74 3.90
                 4.74 2.34 4.60 2.34 4.60 2.02 4.84 2.02 4.84 1.46 5.87 1.46 ;
        POLYGON  3.64 2.96 1.88 2.96 1.88 3.90 1.56 3.90 1.56 2.64 2.50 2.64
                 2.50 1.22 2.82 1.22 2.82 2.64 3.64 2.64 ;
        RECT  1.12 1.22 2.14 1.54 ;
    END
END tbufh_1

MACRO tbufh_0
    CLASS CORE ;
    FOREIGN tbufh_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.32 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.23  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.29 4.54 0.80 4.54 0.80 3.10 1.24 3.10 1.24 4.22 6.97 4.22
                 6.97 2.66 6.86 2.66 6.86 2.34 7.29 2.34 ;
        END
    END a
    PIN en
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.02  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.12 2.40 1.06 2.40 1.06 2.72 0.74 2.72 0.74 2.08 1.12 2.08 ;
        END
    END en
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.35  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.49 1.54 4.37 1.54 4.28 1.63 4.28 2.72 4.32 2.72 4.32 3.90
                 3.77 3.90 3.77 3.58 4.00 3.58 4.00 3.04 3.96 3.04 3.96 2.40
                 3.94 2.40 3.94 2.08 3.96 2.08 3.96 1.43 4.17 1.22 4.49 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 0.90 7.38 0.90 7.38 1.14 7.06 1.14 7.06 0.90 6.66 0.90
                 6.66 1.14 6.34 1.14 6.34 0.90 5.17 0.90 5.17 1.14 4.85 1.14
                 4.85 0.90 3.79 0.90 3.79 1.14 3.47 1.14 3.47 0.90 0.74 0.90
                 0.74 1.58 0.42 1.58 0.42 0.90 0.00 0.90 0.00 -0.90 8.32 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 8.32 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  8.08 4.34 7.76 4.34 7.76 1.78 6.51 1.78 6.51 2.65 5.48 2.65
                 5.48 2.33 6.19 2.33 6.19 1.46 7.76 1.46 7.76 1.22 8.08 1.22 ;
        RECT  5.44 3.58 6.44 3.90 ;
        POLYGON  5.87 1.78 5.16 1.78 5.16 2.34 5.06 2.34 5.06 3.90 4.74 3.90
                 4.74 2.34 4.60 2.34 4.60 2.02 4.84 2.02 4.84 1.46 5.87 1.46 ;
        POLYGON  3.64 2.96 1.88 2.96 1.88 3.90 1.56 3.90 1.56 2.64 2.50 2.64
                 2.50 1.22 2.82 1.22 2.82 2.64 3.64 2.64 ;
        RECT  1.12 1.22 2.14 1.54 ;
    END
END tbufh_0

MACRO sdffpsqb_4
    CLASS CORE ;
    FOREIGN sdffpsqb_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.04 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  12.76 2.68 13.72 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.62 4.32 3.04 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  22.88 3.04 22.84 3.04 22.84 4.54 21.12 4.54 21.12 4.22
                 22.52 4.22 22.52 2.72 22.56 2.72 22.56 1.84 21.12 1.84
                 21.12 1.52 22.88 1.52 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.02  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.92 2.52 8.06 2.52 8.06 2.20 8.48 2.20 8.48 2.08 8.92 2.08 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.80 1.12 2.44 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  23.04 0.90 22.14 0.90 22.14 1.20 21.82 1.20 21.82 0.90
                 18.68 0.90 18.68 1.54 18.36 1.54 18.36 0.90 12.18 0.90
                 12.18 1.48 11.86 1.48 11.86 0.90 1.31 0.90 1.31 1.12 0.99 1.12
                 0.99 0.90 0.00 0.90 0.00 -0.90 23.04 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  23.04 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.22 1.32 4.22
                 1.32 4.86 11.86 4.86 11.86 4.16 12.18 4.16 12.18 4.86
                 14.02 4.86 14.02 4.64 14.34 4.64 14.34 4.86 17.66 4.86
                 17.66 4.62 17.98 4.62 17.98 4.86 19.74 4.86 19.74 4.00
                 20.06 4.00 20.06 4.86 23.04 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  22.14 2.48 20.76 2.48 20.76 4.54 20.44 4.54 20.44 3.12
                 19.36 3.12 19.36 4.54 19.04 4.54 19.04 3.12 18.18 3.12
                 18.18 2.80 20.44 2.80 20.44 1.52 20.76 1.52 20.76 2.16
                 22.14 2.16 ;
        POLYGON  20.12 2.48 17.86 2.48 17.86 3.64 16.50 3.64 16.50 4.48
                 16.18 4.48 16.18 3.32 17.54 3.32 17.54 2.48 16.18 2.48
                 16.18 1.22 16.50 1.22 16.50 2.16 20.12 2.16 ;
        RECT  19.06 1.22 20.06 1.54 ;
        POLYGON  18.68 4.54 18.36 4.54 18.36 4.28 17.20 4.28 17.20 4.48
                 16.88 4.48 16.88 3.96 18.36 3.96 18.36 3.58 18.68 3.58 ;
        RECT  16.88 1.22 17.98 1.54 ;
        POLYGON  15.80 1.54 13.56 1.54 13.56 2.18 13.24 2.18 13.24 1.22
                 15.80 1.22 ;
        RECT  13.24 4.00 15.80 4.32 ;
        POLYGON  15.76 3.68 14.80 3.68 14.80 3.36 15.44 3.36 15.44 2.18
                 14.80 2.18 14.80 1.86 15.76 1.86 ;
        POLYGON  14.56 2.92 14.36 2.92 14.36 3.68 12.88 3.68 12.88 4.32
                 12.56 4.32 12.56 3.68 12.12 3.68 12.12 2.90 10.38 2.90
                 10.38 3.01 10.06 3.01 10.06 2.58 12.12 2.58 12.12 1.80
                 12.56 1.80 12.56 1.58 12.88 1.58 12.88 2.12 12.44 2.12
                 12.44 3.36 14.04 3.36 14.04 2.58 14.56 2.58 ;
        RECT  10.48 1.24 11.48 1.56 ;
        RECT  10.02 3.47 11.48 3.79 ;
        POLYGON  10.98 4.54 8.68 4.54 8.68 3.90 5.96 3.90 5.96 1.86 6.28 1.86
                 6.28 3.58 9.00 3.58 9.00 4.22 10.98 4.22 ;
        POLYGON  10.10 2.18 9.64 2.18 9.64 3.90 9.32 3.90 9.32 3.16 6.60 3.16
                 6.60 2.70 6.92 2.70 6.92 2.84 9.32 2.84 9.32 1.86 9.78 1.86
                 9.78 1.22 10.10 1.22 ;
        RECT  4.58 1.22 9.40 1.54 ;
        RECT  4.58 4.22 8.36 4.54 ;
        RECT  6.66 1.86 7.66 2.18 ;
        POLYGON  5.60 2.18 1.82 2.18 1.82 1.22 2.14 1.22 2.14 1.86 5.60 1.86 ;
        RECT  2.50 3.58 5.60 3.90 ;
        RECT  2.50 1.22 4.20 1.54 ;
        POLYGON  4.20 4.54 1.82 4.54 1.82 3.58 2.14 3.58 2.14 4.22 4.20 4.22 ;
        POLYGON  3.00 3.08 0.48 3.08 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.76 2.68 2.76
                 2.68 2.62 3.00 2.62 ;
    END
END sdffpsqb_4

MACRO sdffpsqb_2
    CLASS CORE ;
    FOREIGN sdffpsqb_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  12.76 2.68 13.72 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.62 4.32 3.04 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.81  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  22.24 3.04 22.18 3.04 22.18 4.54 21.86 4.54 21.86 1.25
                 22.18 1.25 22.18 2.72 22.24 2.72 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.02  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.92 2.52 8.06 2.52 8.06 2.20 8.48 2.20 8.48 2.08 8.92 2.08 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.80 1.12 2.44 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  22.40 0.90 21.44 0.90 21.44 1.43 21.12 1.43 21.12 0.90
                 18.68 0.90 18.68 1.54 18.36 1.54 18.36 0.90 12.18 0.90
                 12.18 1.48 11.86 1.48 11.86 0.90 1.29 0.90 1.29 1.12 0.97 1.12
                 0.97 0.90 0.00 0.90 0.00 -0.90 22.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  22.40 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.22 1.32 4.22
                 1.32 4.86 11.86 4.86 11.86 4.16 12.18 4.16 12.18 4.86
                 14.02 4.86 14.02 4.64 14.34 4.64 14.34 4.86 17.66 4.86
                 17.66 4.62 17.98 4.62 17.98 4.86 19.74 4.86 19.74 4.22
                 20.06 4.22 20.06 4.86 22.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  21.54 2.99 20.76 2.99 20.76 4.54 20.44 4.54 20.44 3.12
                 19.36 3.12 19.36 4.54 19.04 4.54 19.04 3.12 18.18 3.12
                 18.18 2.80 20.44 2.80 20.44 1.52 20.76 1.52 20.76 2.66
                 21.54 2.66 ;
        POLYGON  20.08 2.48 17.86 2.48 17.86 3.64 16.50 3.64 16.50 4.48
                 16.18 4.48 16.18 3.32 17.54 3.32 17.54 2.48 16.18 2.48
                 16.18 1.22 16.50 1.22 16.50 2.16 20.08 2.16 ;
        RECT  19.06 1.22 20.06 1.54 ;
        POLYGON  18.68 4.54 18.36 4.54 18.36 4.28 17.20 4.28 17.20 4.48
                 16.88 4.48 16.88 3.96 18.36 3.96 18.36 3.58 18.68 3.58 ;
        RECT  16.88 1.22 17.98 1.54 ;
        POLYGON  15.80 1.54 13.56 1.54 13.56 2.18 13.24 2.18 13.24 1.22
                 15.80 1.22 ;
        RECT  13.24 4.00 15.80 4.32 ;
        POLYGON  15.76 3.68 14.80 3.68 14.80 3.36 15.44 3.36 15.44 2.18
                 14.80 2.18 14.80 1.86 15.76 1.86 ;
        POLYGON  14.56 2.92 14.36 2.92 14.36 3.68 12.88 3.68 12.88 4.32
                 12.56 4.32 12.56 3.68 12.12 3.68 12.12 2.90 10.38 2.90
                 10.38 3.01 10.06 3.01 10.06 2.58 12.12 2.58 12.12 1.80
                 12.56 1.80 12.56 1.58 12.88 1.58 12.88 2.12 12.44 2.12
                 12.44 3.36 14.04 3.36 14.04 2.58 14.56 2.58 ;
        RECT  10.48 1.24 11.48 1.56 ;
        RECT  10.02 3.58 11.48 3.90 ;
        POLYGON  10.98 4.54 8.68 4.54 8.68 3.90 5.96 3.90 5.96 1.86 6.28 1.86
                 6.28 3.58 9.00 3.58 9.00 4.22 10.98 4.22 ;
        POLYGON  10.10 2.18 9.64 2.18 9.64 3.90 9.32 3.90 9.32 3.16 6.60 3.16
                 6.60 2.70 6.92 2.70 6.92 2.84 9.32 2.84 9.32 1.86 9.78 1.86
                 9.78 1.22 10.10 1.22 ;
        RECT  4.58 1.22 9.40 1.54 ;
        RECT  4.58 4.22 8.36 4.54 ;
        RECT  6.66 1.86 7.66 2.18 ;
        POLYGON  5.60 2.18 1.82 2.18 1.82 1.22 2.14 1.22 2.14 1.86 5.60 1.86 ;
        RECT  2.50 3.58 5.60 3.90 ;
        RECT  2.50 1.22 4.20 1.54 ;
        POLYGON  4.20 4.54 1.82 4.54 1.82 3.58 2.14 3.58 2.14 4.22 4.20 4.22 ;
        POLYGON  3.00 3.08 0.48 3.08 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.76 2.68 2.76
                 2.68 2.62 3.00 2.62 ;
    END
END sdffpsqb_2

MACRO sdffpsqb_1
    CLASS CORE ;
    FOREIGN sdffpsqb_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  12.76 2.68 13.72 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.62 4.32 3.04 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.31  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  22.24 3.04 22.18 3.04 22.18 4.54 21.86 4.54 21.86 1.52
                 22.18 1.52 22.18 2.72 22.24 2.72 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.02  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.92 2.52 8.06 2.52 8.06 2.20 8.48 2.20 8.48 2.08 8.92 2.08 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.80 1.12 2.44 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  22.40 0.90 21.44 0.90 21.44 1.54 21.12 1.54 21.12 0.90
                 18.68 0.90 18.68 1.54 18.36 1.54 18.36 0.90 12.18 0.90
                 12.18 1.48 11.86 1.48 11.86 0.90 1.29 0.90 1.29 1.12 0.97 1.12
                 0.97 0.90 0.00 0.90 0.00 -0.90 22.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  22.40 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.22 1.32 4.22
                 1.32 4.86 11.86 4.86 11.86 4.16 12.18 4.16 12.18 4.86
                 14.02 4.86 14.02 4.64 14.34 4.64 14.34 4.86 17.66 4.86
                 17.66 4.62 17.98 4.62 17.98 4.86 19.74 4.86 19.74 4.22
                 20.06 4.22 20.06 4.86 22.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  21.54 4.54 20.44 4.54 20.44 3.12 19.36 3.12 19.36 4.54
                 19.04 4.54 19.04 3.12 18.18 3.12 18.18 2.80 20.44 2.80
                 20.44 1.52 20.76 1.52 20.76 4.22 21.22 4.22 21.22 2.66
                 21.54 2.66 ;
        POLYGON  20.08 2.48 17.86 2.48 17.86 3.64 16.50 3.64 16.50 4.48
                 16.18 4.48 16.18 3.32 17.54 3.32 17.54 2.48 16.18 2.48
                 16.18 1.22 16.50 1.22 16.50 2.16 20.08 2.16 ;
        RECT  19.06 1.22 20.06 1.54 ;
        POLYGON  18.68 4.54 18.36 4.54 18.36 4.28 17.20 4.28 17.20 4.48
                 16.88 4.48 16.88 3.96 18.36 3.96 18.36 3.58 18.68 3.58 ;
        RECT  16.88 1.22 17.98 1.54 ;
        POLYGON  15.80 1.54 13.56 1.54 13.56 2.18 13.24 2.18 13.24 1.22
                 15.80 1.22 ;
        RECT  13.24 4.00 15.80 4.32 ;
        POLYGON  15.76 3.68 14.80 3.68 14.80 3.36 15.44 3.36 15.44 2.18
                 14.80 2.18 14.80 1.86 15.76 1.86 ;
        POLYGON  14.56 2.92 14.36 2.92 14.36 3.68 12.88 3.68 12.88 4.32
                 12.56 4.32 12.56 3.68 12.12 3.68 12.12 2.90 10.38 2.90
                 10.38 3.01 10.06 3.01 10.06 2.58 12.12 2.58 12.12 1.80
                 12.56 1.80 12.56 1.58 12.88 1.58 12.88 2.12 12.44 2.12
                 12.44 3.36 14.04 3.36 14.04 2.58 14.56 2.58 ;
        RECT  10.48 1.24 11.48 1.56 ;
        RECT  10.02 3.58 11.48 3.90 ;
        POLYGON  10.98 4.54 8.68 4.54 8.68 3.90 5.96 3.90 5.96 1.86 6.28 1.86
                 6.28 3.58 9.00 3.58 9.00 4.22 10.98 4.22 ;
        POLYGON  10.10 2.18 9.64 2.18 9.64 3.90 9.32 3.90 9.32 3.16 6.60 3.16
                 6.60 2.70 6.92 2.70 6.92 2.84 9.32 2.84 9.32 1.86 9.78 1.86
                 9.78 1.22 10.10 1.22 ;
        RECT  4.58 1.22 9.40 1.54 ;
        RECT  4.58 4.22 8.36 4.54 ;
        RECT  6.66 1.86 7.66 2.18 ;
        POLYGON  5.60 2.18 1.82 2.18 1.82 1.22 2.14 1.22 2.14 1.86 5.60 1.86 ;
        RECT  2.50 3.58 5.60 3.90 ;
        RECT  2.50 1.22 4.20 1.54 ;
        POLYGON  4.20 4.54 1.82 4.54 1.82 3.58 2.14 3.58 2.14 4.22 4.20 4.22 ;
        POLYGON  3.00 3.08 0.48 3.08 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.76 2.68 2.76
                 2.68 2.62 3.00 2.62 ;
    END
END sdffpsqb_1

MACRO sdffpsq_4
    CLASS CORE ;
    FOREIGN sdffpsq_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.04 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  12.76 2.68 13.72 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.62 4.32 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  22.84 4.54 22.52 4.54 22.52 3.04 21.44 3.04 21.44 4.54
                 21.12 4.54 21.12 1.22 21.44 1.22 21.44 2.72 22.52 2.72
                 22.52 1.22 22.84 1.22 ;
        END
    END q
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.02  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.92 2.52 8.06 2.52 8.06 2.20 8.48 2.20 8.48 2.08 8.92 2.08 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.80 1.12 2.44 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  23.04 0.90 22.14 0.90 22.14 1.54 21.82 1.54 21.82 0.90
                 18.68 0.90 18.68 1.54 18.36 1.54 18.36 0.90 12.18 0.90
                 12.18 1.48 11.86 1.48 11.86 0.90 1.31 0.90 1.31 1.12 0.99 1.12
                 0.99 0.90 0.00 0.90 0.00 -0.90 23.04 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  23.04 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.22 1.32 4.22
                 1.32 4.86 11.86 4.86 11.86 4.16 12.18 4.16 12.18 4.86
                 14.02 4.86 14.02 4.64 14.34 4.64 14.34 4.86 17.66 4.86
                 17.66 4.62 17.98 4.62 17.98 4.86 19.74 4.86 19.74 4.00
                 20.06 4.00 20.06 4.86 21.82 4.86 21.82 3.58 22.14 3.58
                 22.14 4.86 23.04 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.76 4.54 20.44 4.54 20.44 3.12 19.36 3.12 19.36 4.54
                 19.04 4.54 19.04 3.12 18.18 3.12 18.18 2.80 20.44 2.80
                 20.44 1.22 20.76 1.22 ;
        POLYGON  20.12 2.48 17.86 2.48 17.86 3.64 16.50 3.64 16.50 4.48
                 16.18 4.48 16.18 3.32 17.54 3.32 17.54 2.48 16.18 2.48
                 16.18 1.22 16.50 1.22 16.50 2.16 20.12 2.16 ;
        RECT  19.06 1.22 20.06 1.54 ;
        POLYGON  18.68 4.54 18.36 4.54 18.36 4.28 17.20 4.28 17.20 4.48
                 16.88 4.48 16.88 3.96 18.36 3.96 18.36 3.58 18.68 3.58 ;
        RECT  16.88 1.22 17.98 1.54 ;
        RECT  13.24 1.22 15.80 1.54 ;
        RECT  13.24 4.00 15.80 4.32 ;
        POLYGON  15.76 3.68 14.80 3.68 14.80 3.36 15.44 3.36 15.44 2.18
                 14.80 2.18 14.80 1.86 15.76 1.86 ;
        POLYGON  14.56 2.92 14.36 2.92 14.36 3.68 12.88 3.68 12.88 4.32
                 12.56 4.32 12.56 3.68 12.12 3.68 12.12 2.90 10.38 2.90
                 10.38 3.01 10.06 3.01 10.06 2.58 12.12 2.58 12.12 1.80
                 12.56 1.80 12.56 1.58 12.88 1.58 12.88 2.12 12.44 2.12
                 12.44 3.36 14.04 3.36 14.04 2.58 14.56 2.58 ;
        RECT  10.48 1.24 11.48 1.56 ;
        RECT  10.02 3.47 11.48 3.79 ;
        POLYGON  10.98 4.54 8.68 4.54 8.68 3.90 5.96 3.90 5.96 1.86 6.28 1.86
                 6.28 3.58 9.00 3.58 9.00 4.22 10.98 4.22 ;
        POLYGON  10.10 2.18 9.64 2.18 9.64 3.90 9.32 3.90 9.32 3.16 6.60 3.16
                 6.60 2.70 6.92 2.70 6.92 2.84 9.32 2.84 9.32 1.86 9.78 1.86
                 9.78 1.22 10.10 1.22 ;
        RECT  4.58 1.22 9.40 1.54 ;
        RECT  4.58 4.22 8.36 4.54 ;
        RECT  6.66 1.86 7.66 2.18 ;
        POLYGON  5.60 2.18 1.82 2.18 1.82 1.22 2.14 1.22 2.14 1.86 5.60 1.86 ;
        RECT  2.50 3.58 5.60 3.90 ;
        RECT  2.50 1.22 4.20 1.54 ;
        POLYGON  4.20 4.54 1.82 4.54 1.82 3.58 2.14 3.58 2.14 4.22 4.20 4.22 ;
        POLYGON  3.00 3.08 0.48 3.08 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.76 2.68 2.76
                 2.68 2.62 3.00 2.62 ;
    END
END sdffpsq_4

MACRO sdffpsq_2
    CLASS CORE ;
    FOREIGN sdffpsq_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  12.76 2.68 13.72 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.62 4.32 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  22.24 3.04 22.14 3.04 22.14 4.54 21.82 4.54 21.82 1.22
                 22.14 1.22 22.14 2.72 22.24 2.72 ;
        END
    END q
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.02  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.92 2.52 8.06 2.52 8.06 2.20 8.48 2.20 8.48 2.08 8.92 2.08 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.80 1.12 2.44 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  22.40 0.90 21.44 0.90 21.44 1.54 21.12 1.54 21.12 0.90
                 18.68 0.90 18.68 1.54 18.36 1.54 18.36 0.90 12.18 0.90
                 12.18 1.48 11.86 1.48 11.86 0.90 1.31 0.90 1.31 1.12 0.99 1.12
                 0.99 0.90 0.00 0.90 0.00 -0.90 22.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  22.40 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.22 1.32 4.22
                 1.32 4.86 11.86 4.86 11.86 4.16 12.18 4.16 12.18 4.86
                 14.02 4.86 14.02 4.64 14.34 4.64 14.34 4.86 17.66 4.86
                 17.66 4.62 17.98 4.62 17.98 4.86 19.74 4.86 19.74 4.00
                 20.06 4.00 20.06 4.86 21.12 4.86 21.12 3.58 21.44 3.58
                 21.44 4.86 22.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.76 4.54 20.44 4.54 20.44 3.12 19.36 3.12 19.36 4.54
                 19.04 4.54 19.04 3.12 18.18 3.12 18.18 2.80 20.44 2.80
                 20.44 1.22 20.76 1.22 ;
        POLYGON  20.12 2.48 17.86 2.48 17.86 3.64 16.50 3.64 16.50 4.48
                 16.18 4.48 16.18 3.32 17.54 3.32 17.54 2.48 16.18 2.48
                 16.18 1.22 16.50 1.22 16.50 2.16 20.12 2.16 ;
        RECT  19.06 1.22 20.06 1.54 ;
        POLYGON  18.68 4.54 18.36 4.54 18.36 4.28 17.20 4.28 17.20 4.48
                 16.88 4.48 16.88 3.96 18.36 3.96 18.36 3.58 18.68 3.58 ;
        RECT  16.88 1.22 17.98 1.54 ;
        POLYGON  15.80 1.54 13.56 1.54 13.56 2.18 13.24 2.18 13.24 1.22
                 15.80 1.22 ;
        RECT  13.24 4.00 15.80 4.32 ;
        POLYGON  15.76 3.68 14.80 3.68 14.80 3.36 15.44 3.36 15.44 2.18
                 14.80 2.18 14.80 1.86 15.76 1.86 ;
        POLYGON  14.56 2.92 14.36 2.92 14.36 3.68 12.88 3.68 12.88 4.32
                 12.56 4.32 12.56 3.68 12.12 3.68 12.12 2.90 10.38 2.90
                 10.38 3.01 10.06 3.01 10.06 2.58 12.12 2.58 12.12 1.80
                 12.56 1.80 12.56 1.58 12.88 1.58 12.88 2.12 12.44 2.12
                 12.44 3.36 14.04 3.36 14.04 2.58 14.56 2.58 ;
        RECT  10.48 1.24 11.48 1.56 ;
        RECT  10.02 3.47 11.48 3.79 ;
        POLYGON  10.98 4.54 8.68 4.54 8.68 3.90 5.96 3.90 5.96 1.86 6.28 1.86
                 6.28 3.58 9.00 3.58 9.00 4.22 10.98 4.22 ;
        POLYGON  10.10 2.18 9.64 2.18 9.64 3.90 9.32 3.90 9.32 3.16 6.60 3.16
                 6.60 2.70 6.92 2.70 6.92 2.84 9.32 2.84 9.32 1.86 9.78 1.86
                 9.78 1.22 10.10 1.22 ;
        RECT  4.58 1.22 9.40 1.54 ;
        RECT  4.58 4.22 8.36 4.54 ;
        RECT  6.66 1.86 7.66 2.18 ;
        POLYGON  5.60 2.18 1.82 2.18 1.82 1.22 2.14 1.22 2.14 1.86 5.60 1.86 ;
        RECT  2.50 3.58 5.60 3.90 ;
        RECT  2.50 1.22 4.20 1.54 ;
        POLYGON  4.20 4.54 1.82 4.54 1.82 3.58 2.14 3.58 2.14 4.22 4.20 4.22 ;
        POLYGON  3.00 3.08 0.48 3.08 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.76 2.68 2.76
                 2.68 2.62 3.00 2.62 ;
    END
END sdffpsq_2

MACRO sdffpsq_1
    CLASS CORE ;
    FOREIGN sdffpsq_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  12.76 2.68 13.72 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.62 4.32 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  22.24 3.04 22.14 3.04 22.14 4.54 21.82 4.54 21.82 1.22
                 22.14 1.22 22.14 2.72 22.24 2.72 ;
        END
    END q
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.02  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.92 2.52 8.06 2.52 8.06 2.20 8.48 2.20 8.48 2.08 8.92 2.08 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.80 1.12 2.44 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  22.40 0.90 21.44 0.90 21.44 1.54 21.12 1.54 21.12 0.90
                 18.68 0.90 18.68 1.54 18.36 1.54 18.36 0.90 12.18 0.90
                 12.18 1.48 11.86 1.48 11.86 0.90 1.30 0.90 1.30 1.12 0.98 1.12
                 0.98 0.90 0.00 0.90 0.00 -0.90 22.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  22.40 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.22 1.32 4.22
                 1.32 4.86 11.86 4.86 11.86 4.16 12.18 4.16 12.18 4.86
                 14.02 4.86 14.02 4.64 14.34 4.64 14.34 4.86 17.66 4.86
                 17.66 4.62 17.98 4.62 17.98 4.86 19.74 4.86 19.74 4.00
                 20.06 4.00 20.06 4.86 21.12 4.86 21.12 4.22 21.44 4.22
                 21.44 4.86 22.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.76 4.54 20.44 4.54 20.44 3.12 19.36 3.12 19.36 4.54
                 19.04 4.54 19.04 3.12 18.18 3.12 18.18 2.80 20.44 2.80
                 20.44 1.22 20.76 1.22 ;
        POLYGON  20.12 2.48 17.86 2.48 17.86 3.64 16.50 3.64 16.50 4.48
                 16.18 4.48 16.18 3.32 17.54 3.32 17.54 2.48 16.18 2.48
                 16.18 1.22 16.50 1.22 16.50 2.16 20.12 2.16 ;
        RECT  19.06 1.22 20.06 1.54 ;
        POLYGON  18.68 4.54 18.36 4.54 18.36 4.28 17.20 4.28 17.20 4.48
                 16.88 4.48 16.88 3.96 18.36 3.96 18.36 3.58 18.68 3.58 ;
        RECT  16.88 1.22 17.98 1.54 ;
        POLYGON  15.80 1.54 13.56 1.54 13.56 2.18 13.24 2.18 13.24 1.22
                 15.80 1.22 ;
        RECT  13.24 4.00 15.80 4.32 ;
        POLYGON  15.76 3.68 14.80 3.68 14.80 3.36 15.44 3.36 15.44 2.18
                 14.80 2.18 14.80 1.86 15.76 1.86 ;
        POLYGON  14.56 2.92 14.36 2.92 14.36 3.68 12.88 3.68 12.88 4.32
                 12.56 4.32 12.56 3.68 12.12 3.68 12.12 2.90 10.38 2.90
                 10.38 3.01 10.06 3.01 10.06 2.58 12.12 2.58 12.12 1.80
                 12.56 1.80 12.56 1.58 12.88 1.58 12.88 2.12 12.44 2.12
                 12.44 3.36 14.04 3.36 14.04 2.58 14.56 2.58 ;
        RECT  10.48 1.24 11.48 1.56 ;
        RECT  10.02 3.47 11.48 3.79 ;
        POLYGON  10.98 4.54 8.68 4.54 8.68 3.90 5.96 3.90 5.96 1.86 6.28 1.86
                 6.28 3.58 9.00 3.58 9.00 4.22 10.98 4.22 ;
        POLYGON  10.10 2.18 9.64 2.18 9.64 3.90 9.32 3.90 9.32 3.16 6.60 3.16
                 6.60 2.70 6.92 2.70 6.92 2.84 9.32 2.84 9.32 1.86 9.78 1.86
                 9.78 1.22 10.10 1.22 ;
        RECT  4.58 1.22 9.40 1.54 ;
        RECT  4.58 4.22 8.36 4.54 ;
        RECT  6.66 1.86 7.66 2.18 ;
        POLYGON  5.60 2.18 1.82 2.18 1.82 1.22 2.14 1.22 2.14 1.86 5.60 1.86 ;
        RECT  2.50 3.58 5.60 3.90 ;
        RECT  2.50 1.22 4.20 1.54 ;
        POLYGON  4.20 4.54 1.82 4.54 1.82 3.58 2.14 3.58 2.14 4.22 4.20 4.22 ;
        POLYGON  3.00 3.08 0.48 3.08 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.76 2.68 2.76
                 2.68 2.62 3.00 2.62 ;
    END
END sdffpsq_1

MACRO sdffps_4
    CLASS CORE ;
    FOREIGN sdffps_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 25.60 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  12.76 2.68 13.72 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.62 4.32 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  22.84 1.84 21.44 1.84 21.44 2.72 21.60 2.72 21.60 2.94
                 22.84 2.94 22.84 3.26 21.12 3.26 21.12 1.52 22.84 1.52 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  25.44 3.04 24.92 3.04 24.92 4.54 23.20 4.54 23.20 4.22
                 24.60 4.22 24.60 2.72 24.74 2.72 24.74 1.84 23.20 1.84
                 23.20 1.52 25.06 1.52 25.06 2.72 25.44 2.72 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.02  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.92 2.52 8.06 2.52 8.06 2.20 8.48 2.20 8.48 2.08 8.92 2.08 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.80 1.12 2.44 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  25.60 0.90 24.22 0.90 24.22 1.20 23.90 1.20 23.90 0.90
                 22.14 0.90 22.14 1.20 21.82 1.20 21.82 0.90 18.68 0.90
                 18.68 1.54 18.36 1.54 18.36 0.90 12.18 0.90 12.18 1.48
                 11.86 1.48 11.86 0.90 1.31 0.90 1.31 1.12 0.99 1.12 0.99 0.90
                 0.00 0.90 0.00 -0.90 25.60 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  25.60 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.22 1.32 4.22
                 1.32 4.86 11.86 4.86 11.86 4.16 12.18 4.16 12.18 4.86
                 14.02 4.86 14.02 4.64 14.34 4.64 14.34 4.86 17.66 4.86
                 17.66 4.62 17.98 4.62 17.98 4.86 19.74 4.86 19.74 4.00
                 20.06 4.00 20.06 4.86 21.82 4.86 21.82 4.22 22.14 4.22
                 22.14 4.86 25.60 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  24.22 2.48 23.48 2.48 23.48 3.90 20.76 3.90 20.76 4.54
                 20.44 4.54 20.44 3.12 19.36 3.12 19.36 4.54 19.04 4.54
                 19.04 3.12 18.18 3.12 18.18 2.80 20.44 2.80 20.44 1.52
                 20.76 1.52 20.76 3.58 23.16 3.58 23.16 2.16 24.22 2.16 ;
        POLYGON  20.12 2.48 17.86 2.48 17.86 3.64 16.50 3.64 16.50 4.48
                 16.18 4.48 16.18 3.32 17.54 3.32 17.54 2.48 16.18 2.48
                 16.18 1.22 16.50 1.22 16.50 2.16 20.12 2.16 ;
        RECT  19.06 1.22 20.06 1.54 ;
        POLYGON  18.68 4.54 18.36 4.54 18.36 4.28 17.20 4.28 17.20 4.48
                 16.88 4.48 16.88 3.96 18.36 3.96 18.36 3.58 18.68 3.58 ;
        RECT  16.88 1.22 17.98 1.54 ;
        POLYGON  15.80 1.54 13.56 1.54 13.56 2.18 13.24 2.18 13.24 1.22
                 15.80 1.22 ;
        RECT  13.24 4.00 15.80 4.32 ;
        POLYGON  15.76 3.68 14.80 3.68 14.80 3.36 15.44 3.36 15.44 2.18
                 14.80 2.18 14.80 1.86 15.76 1.86 ;
        POLYGON  14.56 2.92 14.36 2.92 14.36 3.68 12.88 3.68 12.88 4.32
                 12.56 4.32 12.56 3.68 12.12 3.68 12.12 2.90 10.38 2.90
                 10.38 3.01 10.06 3.01 10.06 2.58 12.12 2.58 12.12 1.80
                 12.56 1.80 12.56 1.58 12.88 1.58 12.88 2.12 12.44 2.12
                 12.44 3.36 14.04 3.36 14.04 2.58 14.56 2.58 ;
        RECT  10.48 1.24 11.48 1.56 ;
        RECT  10.02 3.47 11.48 3.79 ;
        POLYGON  10.98 4.54 8.68 4.54 8.68 3.90 5.96 3.90 5.96 1.86 6.28 1.86
                 6.28 3.58 9.00 3.58 9.00 4.22 10.98 4.22 ;
        POLYGON  10.10 2.18 9.64 2.18 9.64 3.90 9.32 3.90 9.32 3.16 6.60 3.16
                 6.60 2.70 6.92 2.70 6.92 2.84 9.32 2.84 9.32 1.86 9.78 1.86
                 9.78 1.22 10.10 1.22 ;
        RECT  4.58 1.22 9.40 1.54 ;
        RECT  4.58 4.22 8.36 4.54 ;
        RECT  6.66 1.86 7.66 2.18 ;
        POLYGON  5.60 2.18 1.82 2.18 1.82 1.22 2.14 1.22 2.14 1.86 5.60 1.86 ;
        RECT  2.50 3.58 5.60 3.90 ;
        RECT  2.50 1.22 4.20 1.54 ;
        POLYGON  4.20 4.54 1.82 4.54 1.82 3.58 2.14 3.58 2.14 4.22 4.20 4.22 ;
        POLYGON  3.00 3.08 0.48 3.08 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.76 2.68 2.76
                 2.68 2.62 3.00 2.62 ;
    END
END sdffps_4

MACRO sdffps_2
    CLASS CORE ;
    FOREIGN sdffps_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  12.76 2.68 13.72 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.62 4.32 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.76  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  21.60 2.40 21.44 2.40 21.44 3.26 21.04 3.26 21.04 2.94
                 21.12 2.94 21.12 1.52 21.44 1.52 21.44 2.08 21.60 2.08 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  23.52 3.04 22.94 3.04 22.94 4.54 22.58 4.54 22.58 4.22
                 22.62 4.22 22.62 1.84 22.58 1.84 22.58 1.52 22.94 1.52
                 22.94 2.72 23.52 2.72 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.02  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.92 2.52 8.06 2.52 8.06 2.20 8.48 2.20 8.48 2.08 8.92 2.08 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.80 1.12 2.44 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  23.68 0.90 22.20 0.90 22.20 1.54 21.88 1.54 21.88 0.90
                 18.68 0.90 18.68 1.54 18.36 1.54 18.36 0.90 12.18 0.90
                 12.18 1.48 11.86 1.48 11.86 0.90 1.24 0.90 1.24 1.12 0.92 1.12
                 0.92 0.90 0.00 0.90 0.00 -0.90 23.68 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  23.68 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.22 1.32 4.22
                 1.32 4.86 11.86 4.86 11.86 4.16 12.18 4.16 12.18 4.86
                 14.02 4.86 14.02 4.64 14.34 4.64 14.34 4.86 17.66 4.86
                 17.66 4.62 17.98 4.62 17.98 4.86 19.74 4.86 19.74 4.22
                 20.06 4.22 20.06 4.86 21.85 4.86 21.85 4.22 22.17 4.22
                 22.17 4.86 23.68 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  22.30 3.90 20.76 3.90 20.76 4.54 20.40 4.54 20.40 3.12
                 19.36 3.12 19.36 4.54 19.04 4.54 19.04 3.12 18.18 3.12
                 18.18 2.80 20.40 2.80 20.40 1.52 20.76 1.52 20.76 1.84
                 20.72 1.84 20.72 3.58 21.98 3.58 21.98 2.66 22.30 2.66 ;
        POLYGON  20.08 2.48 17.86 2.48 17.86 3.64 16.50 3.64 16.50 4.48
                 16.18 4.48 16.18 3.32 17.54 3.32 17.54 2.48 16.18 2.48
                 16.18 1.22 16.50 1.22 16.50 2.16 20.08 2.16 ;
        RECT  19.06 1.22 20.06 1.54 ;
        POLYGON  18.68 4.54 18.36 4.54 18.36 4.28 17.20 4.28 17.20 4.48
                 16.88 4.48 16.88 3.96 18.36 3.96 18.36 3.48 18.68 3.48 ;
        RECT  16.88 1.22 17.98 1.54 ;
        POLYGON  15.80 1.54 13.56 1.54 13.56 2.18 13.24 2.18 13.24 1.22
                 15.80 1.22 ;
        RECT  13.24 4.00 15.80 4.32 ;
        POLYGON  15.76 3.68 14.80 3.68 14.80 3.36 15.44 3.36 15.44 2.18
                 14.80 2.18 14.80 1.86 15.76 1.86 ;
        POLYGON  14.56 2.92 14.36 2.92 14.36 3.68 12.88 3.68 12.88 4.32
                 12.56 4.32 12.56 3.68 12.12 3.68 12.12 2.90 10.38 2.90
                 10.38 3.01 10.06 3.01 10.06 2.58 12.12 2.58 12.12 1.80
                 12.56 1.80 12.56 1.58 12.88 1.58 12.88 2.12 12.44 2.12
                 12.44 3.36 14.04 3.36 14.04 2.58 14.56 2.58 ;
        RECT  10.48 1.24 11.48 1.56 ;
        RECT  10.02 3.58 11.48 3.90 ;
        POLYGON  10.98 4.54 8.68 4.54 8.68 3.90 5.96 3.90 5.96 1.86 6.28 1.86
                 6.28 3.58 9.00 3.58 9.00 4.22 10.98 4.22 ;
        POLYGON  10.10 2.18 9.64 2.18 9.64 3.90 9.32 3.90 9.32 3.16 6.60 3.16
                 6.60 2.70 6.92 2.70 6.92 2.84 9.32 2.84 9.32 1.86 9.78 1.86
                 9.78 1.22 10.10 1.22 ;
        RECT  4.58 1.22 9.40 1.54 ;
        RECT  4.58 4.22 8.36 4.54 ;
        RECT  6.66 1.86 7.66 2.18 ;
        POLYGON  5.60 2.18 1.82 2.18 1.82 1.22 2.14 1.22 2.14 1.86 5.60 1.86 ;
        RECT  2.50 3.58 5.60 3.90 ;
        RECT  2.50 1.22 4.20 1.54 ;
        POLYGON  4.20 4.54 1.82 4.54 1.82 3.58 2.14 3.58 2.14 4.22 4.20 4.22 ;
        POLYGON  3.00 3.08 0.48 3.08 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.76 2.68 2.76
                 2.68 2.62 3.00 2.62 ;
    END
END sdffps_2

MACRO sdffps_1
    CLASS CORE ;
    FOREIGN sdffps_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  12.76 2.68 13.72 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.62 4.32 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.28  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  21.60 2.40 21.44 2.40 21.44 3.90 21.12 3.90 21.12 1.52
                 21.44 1.52 21.44 2.08 21.60 2.08 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.40  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  23.52 3.04 22.94 3.04 22.94 4.54 22.62 4.54 22.62 1.52
                 22.94 1.52 22.94 2.72 23.52 2.72 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.02  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.92 2.52 8.06 2.52 8.06 2.20 8.48 2.20 8.48 2.08 8.92 2.08 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.80 1.12 2.44 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  23.68 0.90 22.20 0.90 22.20 1.54 21.88 1.54 21.88 0.90
                 18.68 0.90 18.68 1.54 18.36 1.54 18.36 0.90 12.18 0.90
                 12.18 1.48 11.86 1.48 11.86 0.90 1.29 0.90 1.29 1.12 0.97 1.12
                 0.97 0.90 0.00 0.90 0.00 -0.90 23.68 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  23.68 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.22 1.32 4.22
                 1.32 4.86 11.86 4.86 11.86 4.16 12.18 4.16 12.18 4.86
                 14.02 4.86 14.02 4.64 14.34 4.64 14.34 4.86 17.66 4.86
                 17.66 4.62 17.98 4.62 17.98 4.86 19.74 4.86 19.74 4.22
                 20.06 4.22 20.06 4.86 23.68 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  22.30 4.54 20.44 4.54 20.44 3.12 19.36 3.12 19.36 4.54
                 19.04 4.54 19.04 3.12 18.18 3.12 18.18 2.80 20.44 2.80
                 20.44 1.52 20.76 1.52 20.76 4.22 21.98 4.22 21.98 2.66
                 22.30 2.66 ;
        POLYGON  20.08 2.48 17.86 2.48 17.86 3.64 16.50 3.64 16.50 4.48
                 16.18 4.48 16.18 3.32 17.54 3.32 17.54 2.48 16.18 2.48
                 16.18 1.22 16.50 1.22 16.50 2.16 20.08 2.16 ;
        RECT  19.06 1.22 20.06 1.54 ;
        POLYGON  18.68 4.54 18.36 4.54 18.36 4.28 17.20 4.28 17.20 4.48
                 16.88 4.48 16.88 3.96 18.36 3.96 18.36 3.58 18.68 3.58 ;
        RECT  16.88 1.22 17.98 1.54 ;
        POLYGON  15.80 1.54 13.56 1.54 13.56 2.18 13.24 2.18 13.24 1.22
                 15.80 1.22 ;
        RECT  13.24 4.00 15.80 4.32 ;
        POLYGON  15.76 3.68 14.80 3.68 14.80 3.36 15.44 3.36 15.44 2.18
                 14.80 2.18 14.80 1.86 15.76 1.86 ;
        POLYGON  14.56 2.92 14.36 2.92 14.36 3.68 12.88 3.68 12.88 4.32
                 12.56 4.32 12.56 3.68 12.12 3.68 12.12 2.90 10.38 2.90
                 10.38 3.01 10.06 3.01 10.06 2.58 12.12 2.58 12.12 1.80
                 12.56 1.80 12.56 1.58 12.88 1.58 12.88 2.12 12.44 2.12
                 12.44 3.36 14.04 3.36 14.04 2.58 14.56 2.58 ;
        RECT  10.48 1.24 11.48 1.56 ;
        RECT  10.02 3.58 11.48 3.90 ;
        POLYGON  10.98 4.54 8.68 4.54 8.68 3.90 5.96 3.90 5.96 1.86 6.28 1.86
                 6.28 3.58 9.00 3.58 9.00 4.22 10.98 4.22 ;
        POLYGON  10.10 2.18 9.64 2.18 9.64 3.90 9.32 3.90 9.32 3.16 6.60 3.16
                 6.60 2.70 6.92 2.70 6.92 2.84 9.32 2.84 9.32 1.86 9.78 1.86
                 9.78 1.22 10.10 1.22 ;
        RECT  4.58 1.22 9.40 1.54 ;
        RECT  4.58 4.22 8.36 4.54 ;
        RECT  6.66 1.86 7.66 2.18 ;
        POLYGON  5.60 2.18 1.82 2.18 1.82 1.22 2.14 1.22 2.14 1.86 5.60 1.86 ;
        RECT  2.50 3.58 5.60 3.90 ;
        RECT  2.50 1.22 4.20 1.54 ;
        POLYGON  4.20 4.54 1.82 4.54 1.82 3.58 2.14 3.58 2.14 4.22 4.20 4.22 ;
        POLYGON  3.00 3.08 0.48 3.08 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.76 2.68 2.76
                 2.68 2.62 3.00 2.62 ;
    END
END sdffps_1

MACRO sdffprsqb_4
    CLASS CORE ;
    FOREIGN sdffprsqb_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 28.16 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.96 3.04 15.84 3.04 15.84 2.72 16.64 2.72 16.64 2.50
                 16.96 2.50 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.62 4.56 3.04 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  28.00 4.54 26.26 4.54 26.26 4.22 27.68 4.22 27.68 1.90
                 26.26 1.90 26.26 1.58 28.00 1.58 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.52 3.04 6.80 3.04 6.80 2.60 7.20 2.60 7.20 2.72 7.52 2.72 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  23.16 2.62 23.52 3.26 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.95 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.76 1.12 2.40 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  28.16 0.90 27.28 0.90 27.28 1.23 26.96 1.23 26.96 0.90
                 25.90 0.90 25.90 1.52 25.58 1.52 25.58 0.90 22.94 0.90
                 22.94 1.53 22.62 1.53 22.62 0.90 1.33 0.90 1.33 1.12 1.01 1.12
                 1.01 0.90 0.00 0.90 0.00 -0.90 28.16 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  28.16 6.66 0.00 6.66 0.00 4.86 1.02 4.86 1.02 4.22 1.34 4.22
                 1.34 4.86 3.24 4.86 3.24 4.66 3.56 4.66 3.56 4.86 15.06 4.86
                 15.06 4.14 15.38 4.14 15.38 4.86 17.58 4.86 17.58 4.64
                 17.90 4.64 17.90 4.86 21.14 4.86 21.14 4.60 21.46 4.60
                 21.46 4.86 28.16 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  27.28 3.90 22.84 3.90 22.84 4.54 22.52 4.54 22.52 3.58
                 22.25 3.58 22.25 3.26 22.84 3.26 22.84 3.58 24.88 3.58
                 24.88 1.22 25.20 1.22 25.20 3.58 26.96 3.58 26.96 2.32
                 27.28 2.32 ;
        RECT  23.27 4.22 25.20 4.54 ;
        RECT  23.50 1.22 24.50 1.54 ;
        POLYGON  24.16 2.64 23.84 2.64 23.84 2.24 21.93 2.24 21.93 3.64
                 20.08 3.64 20.08 4.54 19.76 4.54 19.76 3.32 21.61 3.32
                 21.61 2.24 20.19 2.24 20.19 1.28 20.51 1.28 20.51 1.92
                 24.16 1.92 ;
        POLYGON  22.16 4.28 20.78 4.28 20.78 4.44 20.46 4.44 20.46 3.96
                 22.16 3.96 ;
        RECT  20.89 1.28 22.14 1.60 ;
        POLYGON  19.81 1.60 19.49 1.60 19.49 1.54 17.17 1.54 17.17 1.22
                 19.81 1.22 ;
        POLYGON  19.65 2.58 19.13 2.58 19.13 3.00 18.70 3.00 18.70 3.68
                 18.38 3.68 18.38 2.68 18.81 2.68 18.81 2.18 16.45 2.18
                 16.45 1.54 14.62 1.54 14.62 2.40 13.04 2.40 13.04 2.84
                 12.52 2.84 12.52 2.52 12.72 2.52 12.72 2.08 14.30 2.08
                 14.30 1.22 16.77 1.22 16.77 1.86 19.13 1.86 19.13 2.26
                 19.65 2.26 ;
        RECT  16.80 4.00 19.38 4.32 ;
        POLYGON  18.06 3.08 17.88 3.08 17.88 3.68 16.44 3.68 16.44 4.32
                 16.12 4.32 16.12 3.68 15.00 3.68 15.00 3.06 14.12 3.06
                 14.12 2.74 15.00 2.74 15.00 1.86 16.13 1.86 16.13 2.18
                 15.32 2.18 15.32 3.36 17.56 3.36 17.56 2.76 18.06 2.76 ;
        POLYGON  14.68 3.90 13.68 3.90 13.68 3.46 14.00 3.46 14.00 3.58
                 14.68 3.58 ;
        POLYGON  14.16 4.54 11.78 4.54 11.24 4.00 11.24 3.26 8.52 3.26
                 7.74 2.48 7.74 1.86 8.06 1.86 8.06 2.34 8.66 2.94 11.56 2.94
                 11.56 3.86 11.92 4.22 14.16 4.22 ;
        RECT  12.82 1.28 13.98 1.60 ;
        POLYGON  13.30 3.90 12.06 3.90 11.88 3.72 11.88 2.62 9.76 2.62
                 9.76 2.30 11.88 2.30 11.88 1.96 11.98 1.86 12.08 1.86
                 12.08 1.28 12.40 1.28 12.40 2.18 12.20 2.18 12.20 3.58
                 13.30 3.58 ;
        POLYGON  11.70 1.60 11.38 1.60 11.38 1.54 4.62 1.54 4.62 1.22
                 11.70 1.22 ;
        RECT  4.62 4.22 11.00 4.54 ;
        RECT  7.76 3.58 10.32 3.90 ;
        RECT  8.46 1.86 9.46 2.18 ;
        POLYGON  7.26 2.20 6.94 2.20 6.94 2.18 6.32 2.18 6.32 3.90 6.00 3.90
                 6.00 1.86 7.26 1.86 ;
        POLYGON  5.64 2.18 1.86 2.18 1.86 1.22 2.18 1.22 2.18 1.86 5.64 1.86 ;
        POLYGON  5.64 3.72 5.32 3.72 5.32 3.70 2.54 3.70 2.54 3.38 5.64 3.38 ;
        RECT  2.54 1.22 4.24 1.54 ;
        POLYGON  4.24 4.34 1.86 4.34 1.86 3.38 2.18 3.38 2.18 4.02 4.24 4.02 ;
        POLYGON  3.24 3.04 0.48 3.04 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.72 2.92 2.72
                 2.92 2.60 3.24 2.60 ;
    END
END sdffprsqb_4

MACRO sdffprsqb_2
    CLASS CORE ;
    FOREIGN sdffprsqb_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 27.52 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.96 3.04 15.84 3.04 15.84 2.72 16.64 2.72 16.64 2.50
                 16.96 2.50 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.62 4.56 3.04 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.75  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  27.36 2.40 26.88 2.40 26.88 4.54 26.56 4.54 26.56 1.22
                 26.91 1.22 26.91 1.54 26.88 1.54 26.88 2.08 27.36 2.08 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.52 3.04 6.80 3.04 6.80 2.60 7.20 2.60 7.20 2.72 7.52 2.72 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  23.16 2.62 23.52 3.26 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.95 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.76 1.12 2.40 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  27.52 0.90 26.09 0.90 26.09 1.52 25.77 1.52 25.77 0.90
                 23.01 0.90 23.01 1.53 22.69 1.53 22.69 0.90 1.35 0.90
                 1.35 1.12 1.03 1.12 1.03 0.90 0.00 0.90 0.00 -0.90 27.52 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  27.52 6.66 0.00 6.66 0.00 4.86 1.02 4.86 1.02 4.22 1.34 4.22
                 1.34 4.86 3.24 4.86 3.24 4.66 3.56 4.66 3.56 4.86 15.06 4.86
                 15.06 4.14 15.38 4.14 15.38 4.86 17.58 4.86 17.58 4.64
                 17.90 4.64 17.90 4.86 21.14 4.86 21.14 4.60 21.46 4.60
                 21.46 4.86 25.70 4.86 25.70 4.24 26.02 4.24 26.02 4.86
                 27.52 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  26.13 2.57 25.27 2.57 25.27 3.90 22.84 3.90 22.84 4.54
                 22.52 4.54 22.52 3.58 22.25 3.58 22.25 3.26 22.84 3.26
                 22.84 3.58 24.95 3.58 24.95 1.22 25.27 1.22 25.27 2.25
                 26.13 2.25 ;
        RECT  23.27 4.22 25.20 4.54 ;
        RECT  23.57 1.22 24.57 1.54 ;
        POLYGON  24.16 2.64 23.84 2.64 23.84 2.24 21.93 2.24 21.93 3.64
                 20.08 3.64 20.08 4.54 19.76 4.54 19.76 3.32 21.61 3.32
                 21.61 2.24 20.19 2.24 20.19 1.28 20.51 1.28 20.51 1.92
                 24.16 1.92 ;
        RECT  20.89 1.28 22.21 1.60 ;
        POLYGON  22.16 4.28 20.78 4.28 20.78 4.44 20.46 4.44 20.46 3.96
                 22.16 3.96 ;
        POLYGON  19.81 1.60 19.49 1.60 19.49 1.54 17.17 1.54 17.17 1.22
                 19.81 1.22 ;
        POLYGON  19.65 2.58 19.13 2.58 19.13 3.00 18.70 3.00 18.70 3.68
                 18.38 3.68 18.38 2.68 18.81 2.68 18.81 2.18 16.45 2.18
                 16.45 1.54 14.62 1.54 14.62 2.40 13.04 2.40 13.04 2.84
                 12.52 2.84 12.52 2.52 12.72 2.52 12.72 2.08 14.30 2.08
                 14.30 1.22 16.77 1.22 16.77 1.86 19.13 1.86 19.13 2.26
                 19.65 2.26 ;
        RECT  16.80 4.00 19.38 4.32 ;
        POLYGON  18.06 3.08 17.88 3.08 17.88 3.68 16.44 3.68 16.44 4.32
                 16.12 4.32 16.12 3.68 15.00 3.68 15.00 3.06 14.12 3.06
                 14.12 2.74 15.00 2.74 15.00 1.86 16.13 1.86 16.13 2.18
                 15.32 2.18 15.32 3.36 17.56 3.36 17.56 2.76 18.06 2.76 ;
        POLYGON  14.68 3.90 13.68 3.90 13.68 3.46 14.00 3.46 14.00 3.58
                 14.68 3.58 ;
        POLYGON  14.16 4.54 11.78 4.54 11.24 4.00 11.24 3.26 8.52 3.26
                 7.74 2.48 7.74 1.86 8.06 1.86 8.06 2.34 8.66 2.94 11.56 2.94
                 11.56 3.86 11.92 4.22 14.16 4.22 ;
        RECT  12.82 1.28 13.98 1.60 ;
        POLYGON  13.30 3.90 12.06 3.90 11.88 3.72 11.88 2.62 9.76 2.62
                 9.76 2.30 11.88 2.30 11.88 1.96 11.98 1.86 12.08 1.86
                 12.08 1.28 12.40 1.28 12.40 2.18 12.20 2.18 12.20 3.58
                 13.30 3.58 ;
        POLYGON  11.70 1.60 11.38 1.60 11.38 1.54 4.62 1.54 4.62 1.22
                 11.70 1.22 ;
        RECT  4.62 4.22 11.00 4.54 ;
        RECT  7.76 3.58 10.32 3.90 ;
        RECT  8.46 1.86 9.46 2.18 ;
        POLYGON  7.26 2.20 6.94 2.20 6.94 2.18 6.32 2.18 6.32 3.90 6.00 3.90
                 6.00 1.86 7.26 1.86 ;
        POLYGON  5.64 2.18 1.86 2.18 1.86 1.22 2.18 1.22 2.18 1.86 5.64 1.86 ;
        POLYGON  5.64 3.72 5.32 3.72 5.32 3.70 2.54 3.70 2.54 3.38 5.64 3.38 ;
        RECT  2.54 1.22 4.24 1.54 ;
        POLYGON  4.24 4.34 1.86 4.34 1.86 3.38 2.18 3.38 2.18 4.02 4.24 4.02 ;
        POLYGON  3.24 3.04 0.48 3.04 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.72 2.92 2.72
                 2.92 2.60 3.24 2.60 ;
    END
END sdffprsqb_2

MACRO sdffprsqb_1
    CLASS CORE ;
    FOREIGN sdffprsqb_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 27.52 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.96 3.04 15.84 3.04 15.84 2.72 16.64 2.72 16.64 2.50
                 16.96 2.50 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.62 4.56 3.04 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.26  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  27.36 2.40 26.88 2.40 26.88 4.54 26.56 4.54 26.56 1.22
                 26.91 1.22 26.91 1.54 26.88 1.54 26.88 2.08 27.36 2.08 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.52 3.04 6.80 3.04 6.80 2.60 7.20 2.60 7.20 2.72 7.52 2.72 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  23.16 2.62 23.52 3.26 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.95 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.76 1.12 2.40 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  27.52 0.90 26.09 0.90 26.09 1.52 25.77 1.52 25.77 0.90
                 23.01 0.90 23.01 1.53 22.69 1.53 22.69 0.90 1.35 0.90
                 1.35 1.12 1.03 1.12 1.03 0.90 0.00 0.90 0.00 -0.90 27.52 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  27.52 6.66 0.00 6.66 0.00 4.86 1.02 4.86 1.02 4.22 1.34 4.22
                 1.34 4.86 3.24 4.86 3.24 4.66 3.56 4.66 3.56 4.86 15.06 4.86
                 15.06 4.14 15.38 4.14 15.38 4.86 17.58 4.86 17.58 4.64
                 17.90 4.64 17.90 4.86 21.14 4.86 21.14 4.60 21.46 4.60
                 21.46 4.86 25.70 4.86 25.70 4.24 26.02 4.24 26.02 4.86
                 27.52 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  26.13 2.57 25.27 2.57 25.27 3.90 22.84 3.90 22.84 4.54
                 22.52 4.54 22.52 3.58 22.25 3.58 22.25 3.26 22.84 3.26
                 22.84 3.58 24.95 3.58 24.95 1.22 25.27 1.22 25.27 2.25
                 26.13 2.25 ;
        RECT  23.27 4.22 25.20 4.54 ;
        RECT  23.57 1.22 24.57 1.54 ;
        POLYGON  24.16 2.64 23.84 2.64 23.84 2.24 21.93 2.24 21.93 3.64
                 20.08 3.64 20.08 4.54 19.76 4.54 19.76 3.32 21.61 3.32
                 21.61 2.24 20.19 2.24 20.19 1.28 20.51 1.28 20.51 1.92
                 24.16 1.92 ;
        RECT  20.89 1.28 22.21 1.60 ;
        POLYGON  22.16 4.28 20.78 4.28 20.78 4.44 20.46 4.44 20.46 3.96
                 22.16 3.96 ;
        POLYGON  19.81 1.60 19.49 1.60 19.49 1.54 17.17 1.54 17.17 1.22
                 19.81 1.22 ;
        POLYGON  19.65 2.58 19.13 2.58 19.13 3.00 18.70 3.00 18.70 3.68
                 18.38 3.68 18.38 2.68 18.81 2.68 18.81 2.18 16.45 2.18
                 16.45 1.54 14.62 1.54 14.62 2.40 13.04 2.40 13.04 2.84
                 12.52 2.84 12.52 2.52 12.72 2.52 12.72 2.08 14.30 2.08
                 14.30 1.22 16.77 1.22 16.77 1.86 19.13 1.86 19.13 2.26
                 19.65 2.26 ;
        RECT  16.80 4.00 19.38 4.32 ;
        POLYGON  18.06 3.08 17.88 3.08 17.88 3.68 16.44 3.68 16.44 4.32
                 16.12 4.32 16.12 3.68 15.00 3.68 15.00 3.06 14.12 3.06
                 14.12 2.74 15.00 2.74 15.00 1.86 16.13 1.86 16.13 2.18
                 15.32 2.18 15.32 3.36 17.56 3.36 17.56 2.76 18.06 2.76 ;
        POLYGON  14.68 3.90 13.68 3.90 13.68 3.46 14.00 3.46 14.00 3.58
                 14.68 3.58 ;
        POLYGON  14.16 4.54 11.78 4.54 11.24 4.00 11.24 3.26 8.52 3.26
                 7.74 2.48 7.74 1.86 8.06 1.86 8.06 2.34 8.66 2.94 11.56 2.94
                 11.56 3.86 11.92 4.22 14.16 4.22 ;
        RECT  12.82 1.28 13.98 1.60 ;
        POLYGON  13.30 3.90 12.06 3.90 11.88 3.72 11.88 2.62 9.76 2.62
                 9.76 2.30 11.88 2.30 11.88 1.96 11.98 1.86 12.08 1.86
                 12.08 1.28 12.40 1.28 12.40 2.18 12.20 2.18 12.20 3.58
                 13.30 3.58 ;
        POLYGON  11.70 1.60 11.38 1.60 11.38 1.54 4.62 1.54 4.62 1.22
                 11.70 1.22 ;
        RECT  4.62 4.22 11.00 4.54 ;
        RECT  7.76 3.58 10.32 3.90 ;
        RECT  8.46 1.86 9.46 2.18 ;
        POLYGON  7.26 2.20 6.94 2.20 6.94 2.18 6.32 2.18 6.32 3.90 6.00 3.90
                 6.00 1.86 7.26 1.86 ;
        POLYGON  5.64 2.18 1.86 2.18 1.86 1.22 2.18 1.22 2.18 1.86 5.64 1.86 ;
        POLYGON  5.64 3.72 5.32 3.72 5.32 3.70 2.54 3.70 2.54 3.38 5.64 3.38 ;
        RECT  2.54 1.22 4.24 1.54 ;
        POLYGON  4.24 4.34 1.86 4.34 1.86 3.38 2.18 3.38 2.18 4.02 4.24 4.02 ;
        POLYGON  3.24 3.04 0.48 3.04 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.72 2.92 2.72
                 2.92 2.60 3.24 2.60 ;
    END
END sdffprsqb_1

MACRO sdffprsq_4
    CLASS CORE ;
    FOREIGN sdffprsq_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 29.44 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.96 3.04 15.84 3.04 15.84 2.72 16.64 2.72 16.64 2.50
                 16.96 2.50 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.62 4.56 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  28.99 4.54 28.67 4.54 28.67 2.40 27.71 2.40 27.71 3.28
                 27.59 3.28 27.59 4.54 27.27 4.54 27.27 2.96 27.39 2.96
                 27.39 1.54 27.27 1.54 27.27 1.22 27.71 1.22 27.71 2.08
                 28.67 2.08 28.67 1.22 28.99 1.22 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.52 3.04 6.80 3.04 6.80 2.60 7.20 2.60 7.20 2.72 7.52 2.72 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  23.16 2.62 23.52 3.26 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.95 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.76 1.12 2.40 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  29.44 0.90 25.97 0.90 25.97 1.52 25.65 1.52 25.65 0.90
                 23.01 0.90 23.01 1.53 22.69 1.53 22.69 0.90 1.34 0.90
                 1.34 1.12 1.02 1.12 1.02 0.90 0.00 0.90 0.00 -0.90 29.44 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  29.44 6.66 0.00 6.66 0.00 4.86 1.02 4.86 1.02 4.22 1.34 4.22
                 1.34 4.86 3.24 4.86 3.24 4.66 3.56 4.66 3.56 4.86 15.06 4.86
                 15.06 4.14 15.38 4.14 15.38 4.64 17.98 4.64 17.98 4.86
                 21.14 4.86 21.14 4.60 21.46 4.60 21.46 4.86 25.70 4.86
                 25.70 3.58 26.02 3.58 26.02 4.86 27.97 4.86 27.97 3.58
                 28.29 3.58 28.29 4.86 29.44 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  27.07 2.46 26.88 2.46 26.88 4.54 26.56 4.54 26.56 1.22
                 26.91 1.22 26.91 1.54 26.88 1.54 26.88 2.14 27.07 2.14 ;
        POLYGON  26.13 2.57 25.27 2.57 25.27 3.90 22.84 3.90 22.84 4.54
                 22.52 4.54 22.52 3.58 22.25 3.58 22.25 3.26 22.84 3.26
                 22.84 3.58 24.95 3.58 24.95 1.22 25.27 1.22 25.27 2.25
                 26.13 2.25 ;
        RECT  23.27 4.22 25.20 4.54 ;
        RECT  23.57 1.22 24.57 1.54 ;
        POLYGON  24.16 2.64 23.84 2.64 23.84 2.24 21.93 2.24 21.93 3.64
                 20.08 3.64 20.08 4.54 19.76 4.54 19.76 3.32 21.61 3.32
                 21.61 2.24 20.19 2.24 20.19 1.28 20.51 1.28 20.51 1.92
                 24.16 1.92 ;
        RECT  20.89 1.28 22.21 1.60 ;
        POLYGON  22.16 4.28 20.78 4.28 20.78 4.44 20.46 4.44 20.46 3.96
                 22.16 3.96 ;
        POLYGON  19.81 1.60 19.49 1.60 19.49 1.54 17.17 1.54 17.17 1.22
                 19.81 1.22 ;
        POLYGON  19.65 2.58 19.13 2.58 19.13 3.00 18.70 3.00 18.70 3.68
                 18.38 3.68 18.38 2.68 18.81 2.68 18.81 2.18 16.45 2.18
                 16.45 1.54 14.62 1.54 14.62 2.40 13.04 2.40 13.04 2.84
                 12.52 2.84 12.52 2.52 12.72 2.52 12.72 2.08 14.30 2.08
                 14.30 1.22 16.77 1.22 16.77 1.86 19.13 1.86 19.13 2.26
                 19.65 2.26 ;
        RECT  16.80 4.00 19.38 4.32 ;
        POLYGON  18.06 3.08 17.88 3.08 17.88 3.68 16.44 3.68 16.44 4.32
                 16.12 4.32 16.12 3.68 15.00 3.68 15.00 3.06 14.12 3.06
                 14.12 2.74 15.00 2.74 15.00 1.86 16.13 1.86 16.13 2.18
                 15.32 2.18 15.32 3.36 17.56 3.36 17.56 2.76 18.06 2.76 ;
        POLYGON  14.68 3.90 13.68 3.90 13.68 3.46 14.00 3.46 14.00 3.58
                 14.68 3.58 ;
        POLYGON  14.16 4.54 11.78 4.54 11.24 4.00 11.24 3.26 8.52 3.26
                 7.74 2.48 7.74 1.86 8.06 1.86 8.06 2.34 8.66 2.94 11.56 2.94
                 11.56 3.86 11.92 4.22 14.16 4.22 ;
        RECT  12.82 1.28 13.98 1.60 ;
        POLYGON  13.30 3.90 12.06 3.90 11.88 3.72 11.88 2.62 9.76 2.62
                 9.76 2.30 11.88 2.30 11.88 1.96 11.98 1.86 12.08 1.86
                 12.08 1.28 12.40 1.28 12.40 2.18 12.20 2.18 12.20 3.58
                 13.30 3.58 ;
        POLYGON  11.70 1.60 11.38 1.60 11.38 1.54 4.62 1.54 4.62 1.22
                 11.70 1.22 ;
        RECT  4.62 4.22 11.00 4.54 ;
        RECT  7.76 3.58 10.32 3.90 ;
        RECT  8.46 1.86 9.46 2.18 ;
        POLYGON  7.26 2.20 6.94 2.20 6.94 2.18 6.32 2.18 6.32 3.90 6.00 3.90
                 6.00 1.86 7.26 1.86 ;
        POLYGON  5.64 2.18 1.86 2.18 1.86 1.22 2.18 1.22 2.18 1.86 5.64 1.86 ;
        POLYGON  5.64 3.72 5.32 3.72 5.32 3.70 2.54 3.70 2.54 3.38 5.64 3.38 ;
        RECT  2.54 1.22 4.24 1.54 ;
        POLYGON  4.24 4.34 1.86 4.34 1.86 3.38 2.18 3.38 2.18 4.02 4.24 4.02 ;
        POLYGON  3.24 3.04 0.48 3.04 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.72 2.92 2.72
                 2.92 2.60 3.24 2.60 ;
    END
END sdffprsq_4

MACRO sdffprsq_2
    CLASS CORE ;
    FOREIGN sdffprsq_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 28.80 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.96 3.04 15.84 3.04 15.84 2.72 16.64 2.72 16.64 2.50
                 16.96 2.50 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.62 4.56 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  28.00 2.40 27.71 2.40 27.71 3.28 27.59 3.28 27.59 4.21
                 27.27 4.21 27.27 2.96 27.39 2.96 27.39 1.61 27.27 1.61
                 27.27 1.29 27.71 1.29 27.71 2.08 28.00 2.08 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.52 3.04 6.80 3.04 6.80 2.60 7.20 2.60 7.20 2.72 7.52 2.72 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  23.16 2.62 23.52 3.26 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.95 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.76 1.12 2.40 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  28.80 0.90 26.09 0.90 26.09 1.52 25.77 1.52 25.77 0.90
                 23.01 0.90 23.01 1.53 22.69 1.53 22.69 0.90 1.32 0.90
                 1.32 1.12 1.00 1.12 1.00 0.90 0.00 0.90 0.00 -0.90 28.80 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  28.80 6.66 0.00 6.66 0.00 4.86 1.01 4.86 1.01 4.22 1.33 4.22
                 1.33 4.86 3.24 4.86 3.24 4.66 3.56 4.66 3.56 4.86 15.06 4.86
                 15.06 4.14 15.38 4.14 15.38 4.86 17.58 4.86 17.58 4.64
                 17.90 4.64 17.90 4.86 21.14 4.86 21.14 4.60 21.46 4.60
                 21.46 4.86 25.70 4.86 25.70 4.22 26.02 4.22 26.02 4.86
                 27.97 4.86 27.97 3.89 28.29 3.89 28.29 4.86 28.80 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  27.07 2.46 26.88 2.46 26.88 4.54 26.56 4.54 26.56 1.22
                 26.91 1.22 26.91 1.54 26.88 1.54 26.88 2.14 27.07 2.14 ;
        POLYGON  26.13 2.57 25.27 2.57 25.27 3.90 22.84 3.90 22.84 4.54
                 22.52 4.54 22.52 3.58 22.25 3.58 22.25 3.26 22.84 3.26
                 22.84 3.58 24.95 3.58 24.95 1.22 25.27 1.22 25.27 2.25
                 26.13 2.25 ;
        RECT  23.27 4.22 25.20 4.54 ;
        RECT  23.57 1.22 24.57 1.54 ;
        POLYGON  24.16 2.64 23.84 2.64 23.84 2.24 21.93 2.24 21.93 3.64
                 20.08 3.64 20.08 4.54 19.76 4.54 19.76 3.32 21.61 3.32
                 21.61 2.24 20.19 2.24 20.19 1.28 20.51 1.28 20.51 1.92
                 24.16 1.92 ;
        RECT  20.89 1.28 22.21 1.60 ;
        POLYGON  22.16 4.28 20.78 4.28 20.78 4.44 20.46 4.44 20.46 3.96
                 22.16 3.96 ;
        POLYGON  19.81 1.60 19.49 1.60 19.49 1.54 17.17 1.54 17.17 1.22
                 19.81 1.22 ;
        POLYGON  19.65 2.58 19.13 2.58 19.13 3.00 18.70 3.00 18.70 3.68
                 18.38 3.68 18.38 2.68 18.81 2.68 18.81 2.18 16.45 2.18
                 16.45 1.54 14.62 1.54 14.62 2.40 13.04 2.40 13.04 2.84
                 12.52 2.84 12.52 2.52 12.72 2.52 12.72 2.08 14.30 2.08
                 14.30 1.22 16.77 1.22 16.77 1.86 19.13 1.86 19.13 2.26
                 19.65 2.26 ;
        RECT  16.80 4.00 19.38 4.32 ;
        POLYGON  18.06 3.08 17.88 3.08 17.88 3.68 16.44 3.68 16.44 4.32
                 16.12 4.32 16.12 3.68 15.00 3.68 15.00 3.06 14.12 3.06
                 14.12 2.74 15.00 2.74 15.00 1.86 16.13 1.86 16.13 2.18
                 15.32 2.18 15.32 3.36 17.56 3.36 17.56 2.76 18.06 2.76 ;
        POLYGON  14.68 3.90 13.68 3.90 13.68 3.46 14.00 3.46 14.00 3.58
                 14.68 3.58 ;
        POLYGON  14.16 4.54 11.78 4.54 11.24 4.00 11.24 3.26 8.52 3.26
                 7.74 2.48 7.74 1.86 8.06 1.86 8.06 2.34 8.66 2.94 11.56 2.94
                 11.56 3.86 11.92 4.22 14.16 4.22 ;
        RECT  12.82 1.28 13.98 1.60 ;
        POLYGON  13.30 3.90 12.06 3.90 11.88 3.72 11.88 2.62 9.76 2.62
                 9.76 2.30 11.88 2.30 11.88 1.96 11.98 1.86 12.08 1.86
                 12.08 1.28 12.40 1.28 12.40 2.18 12.20 2.18 12.20 3.58
                 13.30 3.58 ;
        POLYGON  11.70 1.60 11.38 1.60 11.38 1.54 4.62 1.54 4.62 1.22
                 11.70 1.22 ;
        RECT  4.62 4.22 11.00 4.54 ;
        RECT  7.76 3.58 10.32 3.90 ;
        RECT  8.46 1.86 9.46 2.18 ;
        POLYGON  7.26 2.20 6.94 2.20 6.94 2.18 6.32 2.18 6.32 3.90 6.00 3.90
                 6.00 1.86 7.26 1.86 ;
        POLYGON  5.64 2.18 1.86 2.18 1.86 1.22 2.18 1.22 2.18 1.86 5.64 1.86 ;
        POLYGON  5.64 3.72 5.32 3.72 5.32 3.70 2.54 3.70 2.54 3.38 5.64 3.38 ;
        RECT  2.54 1.22 4.24 1.54 ;
        POLYGON  4.24 4.34 1.86 4.34 1.86 3.38 2.18 3.38 2.18 4.02 4.24 4.02 ;
        POLYGON  3.24 3.04 0.48 3.04 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.72 2.92 2.72
                 2.92 2.60 3.24 2.60 ;
    END
END sdffprsq_2

MACRO sdffprsq_1
    CLASS CORE ;
    FOREIGN sdffprsq_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 28.80 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.96 3.04 15.84 3.04 15.84 2.72 16.64 2.72 16.64 2.50
                 16.96 2.50 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.62 4.56 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  28.00 2.40 27.71 2.40 27.71 3.28 27.59 3.28 27.59 4.54
                 27.27 4.54 27.27 2.96 27.39 2.96 27.39 1.54 27.27 1.54
                 27.27 1.22 27.71 1.22 27.71 2.08 28.00 2.08 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.52 3.04 6.80 3.04 6.80 2.60 7.20 2.60 7.20 2.72 7.52 2.72 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  23.16 2.62 23.52 3.26 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.95 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.76 1.12 2.40 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  28.80 0.90 26.09 0.90 26.09 1.52 25.77 1.52 25.77 0.90
                 23.01 0.90 23.01 1.53 22.69 1.53 22.69 0.90 1.35 0.90
                 1.35 1.12 1.03 1.12 1.03 0.90 0.00 0.90 0.00 -0.90 28.80 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  28.80 6.66 0.00 6.66 0.00 4.86 1.02 4.86 1.02 4.22 1.34 4.22
                 1.34 4.86 3.24 4.86 3.24 4.66 3.56 4.66 3.56 4.86 15.06 4.86
                 15.06 4.14 15.38 4.14 15.38 4.86 17.58 4.86 17.58 4.64
                 17.90 4.64 17.90 4.86 21.14 4.86 21.14 4.60 21.46 4.60
                 21.46 4.86 25.70 4.86 25.70 4.24 26.02 4.24 26.02 4.86
                 27.97 4.86 27.97 4.13 28.29 4.13 28.29 4.86 28.80 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  27.07 2.46 26.88 2.46 26.88 4.54 26.56 4.54 26.56 1.22
                 26.91 1.22 26.91 1.54 26.88 1.54 26.88 2.14 27.07 2.14 ;
        POLYGON  26.13 2.57 25.27 2.57 25.27 3.90 22.84 3.90 22.84 4.54
                 22.52 4.54 22.52 3.58 22.25 3.58 22.25 3.26 22.84 3.26
                 22.84 3.58 24.95 3.58 24.95 1.22 25.27 1.22 25.27 2.25
                 26.13 2.25 ;
        RECT  23.27 4.22 25.20 4.54 ;
        RECT  23.57 1.22 24.57 1.54 ;
        POLYGON  24.16 2.64 23.84 2.64 23.84 2.24 21.93 2.24 21.93 3.64
                 20.08 3.64 20.08 4.54 19.76 4.54 19.76 3.32 21.61 3.32
                 21.61 2.24 20.19 2.24 20.19 1.28 20.51 1.28 20.51 1.92
                 24.16 1.92 ;
        RECT  20.89 1.28 22.21 1.60 ;
        POLYGON  22.16 4.28 20.78 4.28 20.78 4.44 20.46 4.44 20.46 3.96
                 22.16 3.96 ;
        POLYGON  19.81 1.60 19.49 1.60 19.49 1.54 17.17 1.54 17.17 1.22
                 19.81 1.22 ;
        POLYGON  19.65 2.58 19.13 2.58 19.13 3.00 18.70 3.00 18.70 3.68
                 18.38 3.68 18.38 2.68 18.81 2.68 18.81 2.18 16.45 2.18
                 16.45 1.54 14.62 1.54 14.62 2.40 13.04 2.40 13.04 2.84
                 12.52 2.84 12.52 2.52 12.72 2.52 12.72 2.08 14.30 2.08
                 14.30 1.22 16.77 1.22 16.77 1.86 19.13 1.86 19.13 2.26
                 19.65 2.26 ;
        RECT  16.80 4.00 19.38 4.32 ;
        POLYGON  18.06 3.08 17.88 3.08 17.88 3.68 16.44 3.68 16.44 4.32
                 16.12 4.32 16.12 3.68 15.00 3.68 15.00 3.06 14.12 3.06
                 14.12 2.74 15.00 2.74 15.00 1.86 16.13 1.86 16.13 2.18
                 15.32 2.18 15.32 3.36 17.56 3.36 17.56 2.76 18.06 2.76 ;
        POLYGON  14.68 3.90 13.68 3.90 13.68 3.46 14.00 3.46 14.00 3.58
                 14.68 3.58 ;
        POLYGON  14.16 4.54 11.78 4.54 11.24 4.00 11.24 3.26 8.52 3.26
                 7.74 2.48 7.74 1.86 8.06 1.86 8.06 2.34 8.66 2.94 11.56 2.94
                 11.56 3.86 11.92 4.22 14.16 4.22 ;
        RECT  12.82 1.28 13.98 1.60 ;
        POLYGON  13.30 3.90 12.06 3.90 11.88 3.72 11.88 2.62 9.76 2.62
                 9.76 2.30 11.88 2.30 11.88 1.96 11.98 1.86 12.08 1.86
                 12.08 1.28 12.40 1.28 12.40 2.18 12.20 2.18 12.20 3.58
                 13.30 3.58 ;
        POLYGON  11.70 1.60 11.38 1.60 11.38 1.54 4.62 1.54 4.62 1.22
                 11.70 1.22 ;
        RECT  4.62 4.22 11.00 4.54 ;
        RECT  7.76 3.58 10.32 3.90 ;
        RECT  8.46 1.86 9.46 2.18 ;
        POLYGON  7.26 2.20 6.94 2.20 6.94 2.18 6.32 2.18 6.32 3.90 6.00 3.90
                 6.00 1.86 7.26 1.86 ;
        POLYGON  5.64 2.18 1.86 2.18 1.86 1.22 2.18 1.22 2.18 1.86 5.64 1.86 ;
        POLYGON  5.64 3.72 5.32 3.72 5.32 3.70 2.54 3.70 2.54 3.38 5.64 3.38 ;
        RECT  2.54 1.22 4.24 1.54 ;
        POLYGON  4.24 4.34 1.86 4.34 1.86 3.38 2.18 3.38 2.18 4.02 4.24 4.02 ;
        POLYGON  3.24 3.04 0.48 3.04 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.72 2.92 2.72
                 2.92 2.60 3.24 2.60 ;
    END
END sdffprsq_1

MACRO sdffprs_4
    CLASS CORE ;
    FOREIGN sdffprs_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 32.00 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.96 3.04 15.84 3.04 15.84 2.72 16.64 2.72 16.64 2.50
                 16.96 2.50 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.62 4.56 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  29.52 3.23 27.75 3.23 27.75 2.91 28.96 2.91 28.96 2.72
                 29.20 2.72 29.20 1.96 27.27 1.96 27.27 1.64 29.52 1.64 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  31.84 4.53 29.84 4.53 29.84 4.21 31.52 4.21 31.52 1.90
                 29.84 1.90 29.84 1.58 31.84 1.58 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.52 3.04 6.80 3.04 6.80 2.60 7.20 2.60 7.20 2.72 7.52 2.72 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  23.16 2.62 23.52 3.26 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.95 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.76 1.12 2.40 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  32.00 0.90 30.86 0.90 30.86 1.23 30.54 1.23 30.54 0.90
                 28.29 0.90 28.29 1.23 27.97 1.23 27.97 0.90 25.97 0.90
                 25.97 1.52 25.65 1.52 25.65 0.90 23.01 0.90 23.01 1.53
                 22.69 1.53 22.69 0.90 1.33 0.90 1.33 1.12 1.01 1.12 1.01 0.90
                 0.00 0.90 0.00 -0.90 32.00 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  32.00 6.66 0.00 6.66 0.00 4.86 1.02 4.86 1.02 4.22 1.34 4.22
                 1.34 4.86 3.24 4.86 3.24 4.66 3.56 4.66 3.56 4.86 15.06 4.86
                 15.06 4.14 15.38 4.14 15.38 4.86 17.58 4.86 17.58 4.64
                 17.90 4.64 17.90 4.86 21.14 4.86 21.14 4.60 21.46 4.60
                 21.46 4.86 28.43 4.86 28.43 4.79 28.80 4.79 28.80 4.86
                 32.00 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  30.86 3.88 28.76 3.88 28.76 4.02 25.62 4.02 25.62 3.90
                 22.84 3.90 22.84 4.54 22.52 4.54 22.52 3.58 22.25 3.58
                 22.25 3.26 22.84 3.26 22.84 3.58 24.95 3.58 24.95 1.22
                 25.27 1.22 25.27 2.25 26.13 2.25 26.13 2.57 25.27 2.57
                 25.27 3.58 25.94 3.58 25.94 3.70 28.44 3.70 28.44 3.56
                 30.54 3.56 30.54 2.32 30.86 2.32 ;
        POLYGON  27.07 2.53 26.88 2.53 26.88 3.38 26.56 3.38 26.56 1.22
                 26.91 1.22 26.91 1.54 26.88 1.54 26.88 2.21 27.07 2.21 ;
        RECT  23.27 4.22 25.20 4.54 ;
        RECT  23.57 1.22 24.57 1.54 ;
        POLYGON  24.16 2.64 23.84 2.64 23.84 2.24 21.93 2.24 21.93 3.64
                 20.08 3.64 20.08 4.54 19.76 4.54 19.76 3.32 21.61 3.32
                 21.61 2.24 20.19 2.24 20.19 1.28 20.51 1.28 20.51 1.92
                 24.16 1.92 ;
        RECT  20.89 1.28 22.21 1.60 ;
        POLYGON  22.16 4.28 20.78 4.28 20.78 4.44 20.46 4.44 20.46 3.96
                 22.16 3.96 ;
        POLYGON  19.81 1.60 19.49 1.60 19.49 1.54 17.17 1.54 17.17 1.22
                 19.81 1.22 ;
        POLYGON  19.65 2.58 19.13 2.58 19.13 3.00 18.70 3.00 18.70 3.68
                 18.38 3.68 18.38 2.68 18.81 2.68 18.81 2.18 16.45 2.18
                 16.45 1.54 14.62 1.54 14.62 2.40 13.04 2.40 13.04 2.84
                 12.52 2.84 12.52 2.52 12.72 2.52 12.72 2.08 14.30 2.08
                 14.30 1.22 16.77 1.22 16.77 1.86 19.13 1.86 19.13 2.26
                 19.65 2.26 ;
        RECT  16.80 4.00 19.38 4.32 ;
        POLYGON  18.06 3.08 17.88 3.08 17.88 3.68 16.44 3.68 16.44 4.32
                 16.12 4.32 16.12 3.68 15.00 3.68 15.00 3.06 14.12 3.06
                 14.12 2.74 15.00 2.74 15.00 1.86 16.13 1.86 16.13 2.18
                 15.32 2.18 15.32 3.36 17.56 3.36 17.56 2.76 18.06 2.76 ;
        POLYGON  14.68 3.90 13.68 3.90 13.68 3.46 14.00 3.46 14.00 3.58
                 14.68 3.58 ;
        POLYGON  14.16 4.54 11.78 4.54 11.24 4.00 11.24 3.26 8.52 3.26
                 7.74 2.48 7.74 1.86 8.06 1.86 8.06 2.34 8.66 2.94 11.56 2.94
                 11.56 3.86 11.92 4.22 14.16 4.22 ;
        RECT  12.82 1.28 13.98 1.60 ;
        POLYGON  13.30 3.90 12.06 3.90 11.88 3.72 11.88 2.62 9.76 2.62
                 9.76 2.30 11.88 2.30 11.88 1.96 11.98 1.86 12.08 1.86
                 12.08 1.28 12.40 1.28 12.40 2.18 12.20 2.18 12.20 3.58
                 13.30 3.58 ;
        POLYGON  11.70 1.60 11.38 1.60 11.38 1.54 4.62 1.54 4.62 1.22
                 11.70 1.22 ;
        RECT  4.62 4.22 11.00 4.54 ;
        RECT  7.76 3.58 10.32 3.90 ;
        RECT  8.46 1.86 9.46 2.18 ;
        POLYGON  7.26 2.20 6.94 2.20 6.94 2.18 6.32 2.18 6.32 3.90 6.00 3.90
                 6.00 1.86 7.26 1.86 ;
        POLYGON  5.64 2.18 1.86 2.18 1.86 1.22 2.18 1.22 2.18 1.86 5.64 1.86 ;
        POLYGON  5.64 3.72 5.32 3.72 5.32 3.70 2.54 3.70 2.54 3.38 5.64 3.38 ;
        RECT  2.54 1.22 4.24 1.54 ;
        POLYGON  4.24 4.34 1.86 4.34 1.86 3.38 2.18 3.38 2.18 4.02 4.24 4.02 ;
        POLYGON  3.24 3.04 0.48 3.04 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.72 2.92 2.72
                 2.92 2.60 3.24 2.60 ;
    END
END sdffprs_4

MACRO sdffprs_2
    CLASS CORE ;
    FOREIGN sdffprs_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 29.44 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.96 3.04 15.84 3.04 15.84 2.72 16.64 2.72 16.64 2.50
                 16.96 2.50 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.62 4.56 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  29.28 4.54 28.64 4.54 28.64 4.22 28.96 4.22 28.96 1.54
                 28.64 1.54 28.64 1.22 29.28 1.22 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  28.00 1.76 27.56 1.76 27.56 3.69 27.24 3.69 27.24 1.44
                 28.00 1.44 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.52 3.04 6.80 3.04 6.80 2.60 7.20 2.60 7.20 2.72 7.52 2.72 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  23.16 2.62 23.52 3.26 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.95 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.76 1.12 2.40 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  29.44 0.90 28.26 0.90 28.26 1.12 27.94 1.12 27.94 0.90
                 25.97 0.90 25.97 1.52 25.65 1.52 25.65 0.90 23.01 0.90
                 23.01 1.53 22.69 1.53 22.69 0.90 1.32 0.90 1.32 1.12 1.00 1.12
                 1.00 0.90 0.00 0.90 0.00 -0.90 29.44 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  29.44 6.66 0.00 6.66 0.00 4.86 1.01 4.86 1.01 4.22 1.33 4.22
                 1.33 4.86 3.24 4.86 3.24 4.66 3.56 4.66 3.56 4.86 15.22 4.86
                 15.22 4.14 15.54 4.14 15.54 4.86 17.58 4.86 17.58 4.64
                 17.90 4.64 17.90 4.86 21.14 4.86 21.14 4.60 21.46 4.60
                 21.46 4.86 25.65 4.86 25.65 4.32 25.97 4.32 25.97 4.86
                 29.44 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  28.42 3.98 28.21 3.98 28.21 4.54 26.56 4.54 26.56 1.22
                 26.88 1.22 26.88 4.22 27.89 4.22 27.89 3.66 28.10 3.66
                 28.10 2.14 28.42 2.14 ;
        POLYGON  26.24 2.57 25.27 2.57 25.27 3.90 22.84 3.90 22.84 4.54
                 22.52 4.54 22.52 3.58 22.25 3.58 22.25 3.26 22.84 3.26
                 22.84 3.58 24.95 3.58 24.95 1.22 25.27 1.22 25.27 2.25
                 26.24 2.25 ;
        RECT  23.27 4.22 25.20 4.54 ;
        RECT  23.57 1.22 24.57 1.54 ;
        POLYGON  24.16 2.64 23.84 2.64 23.84 2.24 21.93 2.24 21.93 3.64
                 20.08 3.64 20.08 4.54 19.76 4.54 19.76 3.32 21.61 3.32
                 21.61 2.24 20.19 2.24 20.19 1.28 20.51 1.28 20.51 1.92
                 24.16 1.92 ;
        RECT  20.89 1.28 22.21 1.60 ;
        POLYGON  22.16 4.28 20.78 4.28 20.78 4.44 20.46 4.44 20.46 3.96
                 22.16 3.96 ;
        POLYGON  19.81 1.60 19.49 1.60 19.49 1.54 17.17 1.54 17.17 1.22
                 19.81 1.22 ;
        POLYGON  19.65 2.58 19.13 2.58 19.13 3.00 18.70 3.00 18.70 3.68
                 18.38 3.68 18.38 2.68 18.81 2.68 18.81 2.18 16.45 2.18
                 16.45 1.54 14.62 1.54 14.62 2.40 13.04 2.40 13.04 2.84
                 12.52 2.84 12.52 2.52 12.72 2.52 12.72 2.08 14.30 2.08
                 14.30 1.22 16.77 1.22 16.77 1.86 19.13 1.86 19.13 2.26
                 19.65 2.26 ;
        RECT  16.80 4.00 19.38 4.32 ;
        POLYGON  18.06 3.08 17.88 3.08 17.88 3.68 16.44 3.68 16.44 4.32
                 16.12 4.32 16.12 3.68 15.00 3.68 15.00 3.06 14.12 3.06
                 14.12 2.74 15.00 2.74 15.00 1.86 16.13 1.86 16.13 2.18
                 15.32 2.18 15.32 3.36 17.56 3.36 17.56 2.76 18.06 2.76 ;
        POLYGON  14.68 3.90 13.68 3.90 13.68 3.46 14.00 3.46 14.00 3.58
                 14.68 3.58 ;
        POLYGON  14.16 4.54 11.78 4.54 11.24 4.00 11.24 3.26 8.52 3.26
                 7.74 2.48 7.74 1.86 8.06 1.86 8.06 2.34 8.66 2.94 11.56 2.94
                 11.56 3.86 11.92 4.22 14.16 4.22 ;
        RECT  12.82 1.28 13.98 1.60 ;
        POLYGON  13.30 3.90 12.06 3.90 11.88 3.72 11.88 2.62 9.76 2.62
                 9.76 2.30 11.88 2.30 11.88 1.96 11.98 1.86 12.08 1.86
                 12.08 1.28 12.40 1.28 12.40 2.18 12.20 2.18 12.20 3.58
                 13.30 3.58 ;
        POLYGON  11.70 1.60 11.38 1.60 11.38 1.54 4.62 1.54 4.62 1.22
                 11.70 1.22 ;
        RECT  4.62 4.22 11.00 4.54 ;
        RECT  7.76 3.58 10.32 3.90 ;
        RECT  8.46 1.86 9.46 2.18 ;
        POLYGON  7.26 2.20 6.94 2.20 6.94 2.18 6.32 2.18 6.32 3.90 6.00 3.90
                 6.00 1.86 7.26 1.86 ;
        POLYGON  5.64 2.18 1.86 2.18 1.86 1.22 2.18 1.22 2.18 1.86 5.64 1.86 ;
        POLYGON  5.64 3.72 5.32 3.72 5.32 3.70 2.54 3.70 2.54 3.38 5.64 3.38 ;
        RECT  2.54 1.22 4.24 1.54 ;
        POLYGON  4.24 4.34 1.86 4.34 1.86 3.38 2.18 3.38 2.18 4.02 4.24 4.02 ;
        POLYGON  3.24 3.04 0.48 3.04 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.72 2.92 2.72
                 2.92 2.60 3.24 2.60 ;
    END
END sdffprs_2

MACRO sdffprs_1
    CLASS CORE ;
    FOREIGN sdffprs_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 29.44 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.96 3.04 15.84 3.04 15.84 2.72 16.64 2.72 16.64 2.50
                 16.96 2.50 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.62 4.56 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  28.00 3.04 27.56 3.04 27.56 4.44 27.24 4.44 27.24 1.22
                 27.56 1.22 27.56 2.72 28.00 2.72 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  28.96 4.44 28.64 4.44 28.64 2.40 28.32 2.40 28.32 2.08
                 28.64 2.08 28.64 1.22 28.96 1.22 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.52 3.04 6.80 3.04 6.80 2.60 7.20 2.60 7.20 2.72 7.52 2.72 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  23.16 2.62 23.52 3.26 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.95 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.76 1.12 2.40 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  29.44 0.90 28.26 0.90 28.26 1.34 27.94 1.34 27.94 0.90
                 25.97 0.90 25.97 1.52 25.65 1.52 25.65 0.90 23.01 0.90
                 23.01 1.53 22.69 1.53 22.69 0.90 1.32 0.90 1.32 1.12 1.00 1.12
                 1.00 0.90 0.00 0.90 0.00 -0.90 29.44 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  29.44 6.66 0.00 6.66 0.00 4.86 1.02 4.86 1.02 4.22 1.34 4.22
                 1.34 4.86 3.24 4.86 3.24 4.66 3.56 4.66 3.56 4.86 15.06 4.86
                 15.06 4.14 15.38 4.14 15.38 4.86 17.58 4.86 17.58 4.64
                 17.90 4.64 17.90 4.86 21.14 4.86 21.14 4.60 21.46 4.60
                 21.46 4.86 25.65 4.86 25.65 4.24 25.97 4.24 25.97 4.86
                 27.94 4.86 27.94 4.28 28.26 4.28 28.26 4.86 29.44 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  26.56 1.22 26.88 4.54 ;
        POLYGON  26.13 2.57 25.27 2.57 25.27 3.90 22.84 3.90 22.84 4.54
                 22.52 4.54 22.52 3.58 22.25 3.58 22.25 3.26 22.84 3.26
                 22.84 3.58 24.95 3.58 24.95 1.22 25.27 1.22 25.27 2.25
                 26.13 2.25 ;
        RECT  23.27 4.22 25.20 4.54 ;
        RECT  23.57 1.22 24.57 1.54 ;
        POLYGON  24.16 2.64 23.84 2.64 23.84 2.24 21.93 2.24 21.93 3.64
                 20.08 3.64 20.08 4.54 19.76 4.54 19.76 3.32 21.61 3.32
                 21.61 2.24 20.19 2.24 20.19 1.28 20.51 1.28 20.51 1.92
                 24.16 1.92 ;
        RECT  20.89 1.28 22.21 1.60 ;
        POLYGON  22.16 4.28 20.78 4.28 20.78 4.44 20.46 4.44 20.46 3.96
                 22.16 3.96 ;
        POLYGON  19.81 1.60 19.49 1.60 19.49 1.54 17.17 1.54 17.17 1.22
                 19.81 1.22 ;
        POLYGON  19.65 2.58 19.13 2.58 19.13 3.00 18.70 3.00 18.70 3.68
                 18.38 3.68 18.38 2.68 18.81 2.68 18.81 2.18 16.45 2.18
                 16.45 1.54 14.62 1.54 14.62 2.40 13.04 2.40 13.04 2.84
                 12.52 2.84 12.52 2.52 12.72 2.52 12.72 2.08 14.30 2.08
                 14.30 1.22 16.77 1.22 16.77 1.86 19.13 1.86 19.13 2.26
                 19.65 2.26 ;
        RECT  16.80 4.00 19.38 4.32 ;
        POLYGON  18.06 3.08 17.88 3.08 17.88 3.68 16.44 3.68 16.44 4.32
                 16.12 4.32 16.12 3.68 15.00 3.68 15.00 3.06 14.12 3.06
                 14.12 2.74 15.00 2.74 15.00 1.86 16.13 1.86 16.13 2.18
                 15.32 2.18 15.32 3.36 17.56 3.36 17.56 2.76 18.06 2.76 ;
        POLYGON  14.68 3.90 13.68 3.90 13.68 3.46 14.00 3.46 14.00 3.58
                 14.68 3.58 ;
        POLYGON  14.16 4.54 11.78 4.54 11.24 4.00 11.24 3.26 8.52 3.26
                 7.74 2.48 7.74 1.86 8.06 1.86 8.06 2.34 8.66 2.94 11.56 2.94
                 11.56 3.86 11.92 4.22 14.16 4.22 ;
        RECT  12.82 1.28 13.98 1.60 ;
        POLYGON  13.30 3.90 12.06 3.90 11.88 3.72 11.88 2.62 9.76 2.62
                 9.76 2.30 11.88 2.30 11.88 1.96 11.98 1.86 12.08 1.86
                 12.08 1.28 12.40 1.28 12.40 2.18 12.20 2.18 12.20 3.58
                 13.30 3.58 ;
        POLYGON  11.70 1.60 11.38 1.60 11.38 1.54 4.62 1.54 4.62 1.22
                 11.70 1.22 ;
        RECT  4.62 4.22 11.00 4.54 ;
        RECT  7.76 3.58 10.32 3.90 ;
        RECT  8.46 1.86 9.46 2.18 ;
        POLYGON  7.26 2.20 6.94 2.20 6.94 2.18 6.32 2.18 6.32 3.90 6.00 3.90
                 6.00 1.86 7.26 1.86 ;
        POLYGON  5.64 2.18 1.86 2.18 1.86 1.22 2.18 1.22 2.18 1.86 5.64 1.86 ;
        POLYGON  5.64 3.72 5.32 3.72 5.32 3.70 2.54 3.70 2.54 3.38 5.64 3.38 ;
        RECT  2.54 1.22 4.24 1.54 ;
        POLYGON  4.24 4.34 1.86 4.34 1.86 3.38 2.18 3.38 2.18 4.02 4.24 4.02 ;
        POLYGON  3.24 3.04 0.48 3.04 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.72 2.92 2.72
                 2.92 2.60 3.24 2.60 ;
    END
END sdffprs_1

MACRO sdffprqb_4
    CLASS CORE ;
    FOREIGN sdffprqb_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 26.88 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  13.52 2.72 14.18 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.65 5.28 3.04 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.86  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  26.72 3.04 26.64 3.04 26.64 4.54 24.76 4.54 24.76 4.22
                 26.32 4.22 26.32 1.54 24.76 1.54 24.76 1.22 26.64 1.22
                 26.64 2.72 26.72 2.72 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.44  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  8.48 2.08 8.94 2.62 ;
        END
    END rb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.60 2.65 6.34 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.65 3.04 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  26.88 0.90 23.46 0.90 23.46 1.54 23.14 1.54 23.14 0.90
                 14.04 0.90 14.04 1.14 13.72 1.14 13.72 0.90 1.88 0.90
                 1.88 1.71 0.88 1.71 0.88 0.90 0.00 0.90 0.00 -0.90 26.88 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  26.88 6.66 0.00 6.66 0.00 4.86 21.76 4.86 21.76 4.12
                 22.08 4.12 22.08 4.86 23.26 4.86 23.26 4.56 23.58 4.56
                 23.58 4.86 26.88 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  25.79 2.46 24.40 2.46 24.40 4.08 24.08 4.08 24.08 3.16
                 21.80 3.16 21.80 2.84 24.08 2.84 24.08 1.54 23.84 1.54
                 23.84 1.22 24.40 1.22 24.40 2.14 25.79 2.14 ;
        POLYGON  23.64 2.52 21.48 2.52 21.48 3.48 22.76 3.48 22.76 4.54
                 22.44 4.54 22.44 3.80 20.14 3.80 19.90 4.04 19.90 4.54
                 19.58 4.54 19.58 3.90 20.00 3.48 21.16 3.48 21.16 2.52
                 20.44 2.52 19.68 1.76 19.68 1.22 20.00 1.22 20.00 1.62
                 20.58 2.20 23.64 2.20 ;
        RECT  21.76 1.22 22.76 1.54 ;
        RECT  20.38 1.22 21.38 1.54 ;
        RECT  20.28 4.12 21.38 4.44 ;
        POLYGON  19.74 2.60 19.42 2.60 19.42 3.24 18.76 3.90 17.66 3.90
                 17.66 4.54 13.86 4.54 13.86 4.05 13.71 3.90 12.54 3.90
                 12.54 3.06 11.80 3.06 11.80 2.74 12.86 2.74 12.86 3.58
                 13.85 3.58 14.18 3.91 14.18 4.22 17.34 4.22 17.34 3.58
                 18.62 3.58 19.10 3.10 19.10 2.50 18.78 2.18 16.06 2.18
                 16.06 1.86 18.92 1.86 19.34 2.28 19.74 2.28 ;
        RECT  18.30 1.22 19.30 1.54 ;
        RECT  18.20 4.22 19.20 4.54 ;
        POLYGON  18.78 2.96 17.02 2.96 17.02 3.90 14.50 3.90 14.50 2.18
                 11.48 2.18 11.48 3.26 11.16 3.26 11.16 1.86 14.82 1.86
                 14.82 3.58 16.70 3.58 16.70 2.64 18.78 2.64 ;
        POLYGON  17.92 1.54 15.74 1.54 15.74 2.54 16.28 2.54 16.28 2.86
                 15.42 2.86 15.42 1.22 17.92 1.22 ;
        POLYGON  13.54 4.54 9.88 4.54 9.88 3.90 6.86 3.90 6.86 2.68 7.22 2.32
                 7.22 1.87 7.54 1.87 7.54 2.46 7.18 2.82 7.18 3.58 10.20 3.58
                 10.20 4.22 13.54 4.22 ;
        RECT  12.34 1.22 13.34 1.54 ;
        RECT  11.22 3.58 12.22 3.90 ;
        RECT  10.96 1.22 11.96 1.54 ;
        POLYGON  10.84 3.90 10.52 3.90 10.52 3.26 7.52 3.26 7.52 2.94
                 10.52 2.94 10.52 2.40 10.26 2.40 10.26 1.22 10.58 1.22
                 10.58 2.08 10.84 2.08 ;
        RECT  5.84 1.22 9.88 1.54 ;
        RECT  5.48 4.22 9.56 4.54 ;
        RECT  2.94 1.87 6.86 2.19 ;
        RECT  4.10 3.58 6.50 3.90 ;
        RECT  4.34 1.23 5.34 1.55 ;
        RECT  2.70 4.22 5.10 4.54 ;
        POLYGON  4.26 2.97 3.78 2.97 3.78 3.90 0.18 3.90 0.18 1.87 0.50 1.87
                 0.50 3.58 3.46 3.58 3.46 2.65 4.26 2.65 ;
        RECT  2.26 1.23 3.96 1.55 ;
    END
END sdffprqb_4

MACRO sdffprqb_2
    CLASS CORE ;
    FOREIGN sdffprqb_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 26.24 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  13.52 2.72 14.18 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.65 5.28 3.04 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  26.08 4.13 25.45 4.13 25.45 3.81 25.76 3.81 25.76 1.64
                 25.46 1.64 25.46 1.32 26.08 1.32 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.44  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  8.48 2.08 8.94 2.62 ;
        END
    END rb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.60 2.65 6.34 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.65 3.04 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  26.24 0.90 23.46 0.90 23.46 1.54 23.14 1.54 23.14 0.90
                 14.04 0.90 14.04 1.14 13.72 1.14 13.72 0.90 1.88 0.90
                 1.88 1.71 0.88 1.71 0.88 0.90 0.00 0.90 0.00 -0.90 26.24 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  26.24 6.66 0.00 6.66 0.00 4.86 21.76 4.86 21.76 4.12
                 22.08 4.12 22.08 4.86 23.26 4.86 23.26 4.56 23.58 4.56
                 23.58 4.86 24.76 4.86 24.76 3.79 25.08 3.79 25.08 4.86
                 26.24 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  25.24 2.46 24.36 2.46 24.36 3.76 24.43 3.76 24.43 4.08
                 24.04 4.08 24.04 3.16 21.80 3.16 21.80 2.84 24.04 2.84
                 24.04 1.54 23.84 1.54 23.84 1.22 24.36 1.22 24.36 2.14
                 25.24 2.14 ;
        POLYGON  23.64 2.52 21.48 2.52 21.48 3.48 22.76 3.48 22.76 4.54
                 22.44 4.54 22.44 3.80 20.14 3.80 19.90 4.04 19.90 4.54
                 19.58 4.54 19.58 3.90 20.00 3.48 21.16 3.48 21.16 2.52
                 20.44 2.52 19.68 1.76 19.68 1.22 20.00 1.22 20.00 1.62
                 20.58 2.20 23.64 2.20 ;
        RECT  21.76 1.22 22.76 1.54 ;
        RECT  20.38 1.22 21.38 1.54 ;
        RECT  20.28 4.12 21.38 4.44 ;
        POLYGON  19.74 2.60 19.42 2.60 19.42 3.24 18.76 3.90 17.66 3.90
                 17.66 4.54 13.86 4.54 13.86 4.05 13.71 3.90 12.54 3.90
                 12.54 3.06 11.80 3.06 11.80 2.74 12.86 2.74 12.86 3.58
                 13.85 3.58 14.18 3.91 14.18 4.22 17.34 4.22 17.34 3.58
                 18.62 3.58 19.10 3.10 19.10 2.50 18.78 2.18 16.06 2.18
                 16.06 1.86 18.92 1.86 19.34 2.28 19.74 2.28 ;
        RECT  18.30 1.22 19.30 1.54 ;
        RECT  18.20 4.22 19.20 4.54 ;
        POLYGON  18.78 2.96 17.02 2.96 17.02 3.90 14.50 3.90 14.50 2.18
                 11.48 2.18 11.48 3.26 11.16 3.26 11.16 1.86 14.82 1.86
                 14.82 3.58 16.70 3.58 16.70 2.64 18.78 2.64 ;
        POLYGON  17.92 1.54 15.74 1.54 15.74 2.54 16.28 2.54 16.28 2.86
                 15.42 2.86 15.42 1.22 17.92 1.22 ;
        POLYGON  13.54 4.54 9.88 4.54 9.88 3.90 6.86 3.90 6.86 2.68 7.22 2.32
                 7.22 1.87 7.54 1.87 7.54 2.46 7.18 2.82 7.18 3.58 10.20 3.58
                 10.20 4.22 13.54 4.22 ;
        RECT  12.34 1.22 13.34 1.54 ;
        RECT  11.22 3.58 12.22 3.90 ;
        RECT  10.96 1.22 11.96 1.54 ;
        POLYGON  10.84 3.90 10.52 3.90 10.52 3.26 7.52 3.26 7.52 2.94
                 10.52 2.94 10.52 2.40 10.26 2.40 10.26 1.22 10.58 1.22
                 10.58 2.08 10.84 2.08 ;
        RECT  5.84 1.22 9.88 1.54 ;
        RECT  5.48 4.22 9.56 4.54 ;
        RECT  2.94 1.87 6.86 2.19 ;
        RECT  4.10 3.58 6.50 3.90 ;
        RECT  4.34 1.23 5.34 1.55 ;
        RECT  2.70 4.22 5.10 4.54 ;
        POLYGON  4.26 2.97 3.78 2.97 3.78 3.90 0.18 3.90 0.18 1.87 0.50 1.87
                 0.50 3.58 3.46 3.58 3.46 2.65 4.26 2.65 ;
        RECT  2.26 1.23 3.96 1.55 ;
    END
END sdffprqb_2

MACRO sdffprqb_1
    CLASS CORE ;
    FOREIGN sdffprqb_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 26.24 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  13.52 2.72 14.18 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.65 5.28 3.04 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  26.08 4.06 25.45 4.06 25.45 3.74 25.76 3.74 25.76 1.54
                 25.46 1.54 25.46 1.22 26.08 1.22 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.44  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  8.48 2.08 8.94 2.62 ;
        END
    END rb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.60 2.65 6.34 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.65 3.04 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  26.24 0.90 23.46 0.90 23.46 1.54 23.14 1.54 23.14 0.90
                 14.04 0.90 14.04 1.14 13.72 1.14 13.72 0.90 1.88 0.90
                 1.88 1.71 0.88 1.71 0.88 0.90 0.00 0.90 0.00 -0.90 26.24 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  26.24 6.66 0.00 6.66 0.00 4.86 21.76 4.86 21.76 4.12
                 22.08 4.12 22.08 4.86 23.26 4.86 23.26 4.56 23.58 4.56
                 23.58 4.86 24.76 4.86 24.76 4.56 25.08 4.56 25.08 4.86
                 26.24 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  25.24 2.46 24.36 2.46 24.36 3.76 24.42 3.76 24.42 4.08
                 24.04 4.08 24.04 3.16 21.80 3.16 21.80 2.84 24.04 2.84
                 24.04 1.54 23.84 1.54 23.84 1.22 24.36 1.22 24.36 2.14
                 25.24 2.14 ;
        POLYGON  23.64 2.52 21.48 2.52 21.48 3.48 22.76 3.48 22.76 4.54
                 22.44 4.54 22.44 3.80 20.14 3.80 19.90 4.04 19.90 4.54
                 19.58 4.54 19.58 3.90 20.00 3.48 21.16 3.48 21.16 2.52
                 20.44 2.52 19.68 1.76 19.68 1.22 20.00 1.22 20.00 1.62
                 20.58 2.20 23.64 2.20 ;
        RECT  21.76 1.22 22.76 1.54 ;
        RECT  20.38 1.22 21.38 1.54 ;
        RECT  20.28 4.12 21.38 4.44 ;
        POLYGON  19.74 2.60 19.42 2.60 19.42 3.24 18.76 3.90 17.66 3.90
                 17.66 4.54 13.86 4.54 13.86 4.05 13.71 3.90 12.54 3.90
                 12.54 3.06 11.80 3.06 11.80 2.74 12.86 2.74 12.86 3.58
                 13.85 3.58 14.18 3.91 14.18 4.22 17.34 4.22 17.34 3.58
                 18.62 3.58 19.10 3.10 19.10 2.50 18.78 2.18 16.06 2.18
                 16.06 1.86 18.92 1.86 19.34 2.28 19.74 2.28 ;
        RECT  18.30 1.22 19.30 1.54 ;
        RECT  18.20 4.22 19.20 4.54 ;
        POLYGON  18.78 2.96 17.02 2.96 17.02 3.90 14.50 3.90 14.50 2.18
                 11.48 2.18 11.48 3.26 11.16 3.26 11.16 1.86 14.82 1.86
                 14.82 3.58 16.70 3.58 16.70 2.64 18.78 2.64 ;
        POLYGON  17.92 1.54 15.74 1.54 15.74 2.54 16.28 2.54 16.28 2.86
                 15.42 2.86 15.42 1.22 17.92 1.22 ;
        POLYGON  13.54 4.54 9.88 4.54 9.88 3.90 6.86 3.90 6.86 2.68 7.22 2.32
                 7.22 1.87 7.54 1.87 7.54 2.46 7.18 2.82 7.18 3.58 10.20 3.58
                 10.20 4.22 13.54 4.22 ;
        RECT  12.34 1.22 13.34 1.54 ;
        RECT  11.22 3.58 12.22 3.90 ;
        RECT  10.96 1.22 11.96 1.54 ;
        POLYGON  10.84 3.90 10.52 3.90 10.52 3.26 7.52 3.26 7.52 2.94
                 10.52 2.94 10.52 2.40 10.26 2.40 10.26 1.22 10.58 1.22
                 10.58 2.08 10.84 2.08 ;
        RECT  5.84 1.22 9.88 1.54 ;
        RECT  5.48 4.22 9.56 4.54 ;
        RECT  2.94 1.87 6.86 2.19 ;
        RECT  4.10 3.58 6.50 3.90 ;
        RECT  4.34 1.23 5.34 1.55 ;
        RECT  2.70 4.22 5.10 4.54 ;
        POLYGON  4.26 2.97 3.78 2.97 3.78 3.90 0.18 3.90 0.18 1.87 0.50 1.87
                 0.50 3.58 3.46 3.58 3.46 2.65 4.26 2.65 ;
        RECT  2.26 1.23 3.96 1.55 ;
    END
END sdffprqb_1

MACRO sdffprq_4
    CLASS CORE ;
    FOREIGN sdffprq_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 26.88 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  13.52 2.72 14.18 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.65 5.28 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  26.48 4.54 26.16 4.54 26.16 3.04 25.08 3.04 25.08 4.54
                 24.76 4.54 24.76 1.22 25.08 1.22 25.08 2.72 26.16 2.72
                 26.16 1.22 26.48 1.22 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.44  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  8.48 2.08 8.94 2.62 ;
        END
    END rb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.60 2.65 6.34 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.65 3.04 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  26.88 0.90 25.78 0.90 25.78 1.54 25.46 1.54 25.46 0.90
                 23.46 0.90 23.46 1.54 23.14 1.54 23.14 0.90 14.04 0.90
                 14.04 1.54 13.72 1.54 13.72 0.90 1.88 0.90 1.88 1.71 0.88 1.71
                 0.88 0.90 0.00 0.90 0.00 -0.90 26.88 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  26.88 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 21.76 4.86 21.76 4.22 22.08 4.22 22.08 4.86
                 23.26 4.86 23.26 4.22 23.58 4.22 23.58 4.86 25.46 4.86
                 25.46 3.58 25.78 3.58 25.78 4.86 26.88 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  24.40 4.54 24.08 4.54 24.08 3.16 21.80 3.16 21.80 2.84
                 24.08 2.84 24.08 1.54 23.84 1.54 23.84 1.22 24.40 1.22 ;
        POLYGON  23.64 2.52 21.48 2.52 21.48 3.48 22.76 3.48 22.76 4.54
                 22.44 4.54 22.44 3.80 20.14 3.80 19.90 4.04 19.90 4.54
                 19.58 4.54 19.58 3.90 20.00 3.48 21.16 3.48 21.16 2.52
                 20.44 2.52 19.68 1.76 19.68 1.22 20.00 1.22 20.00 1.62
                 20.58 2.20 23.64 2.20 ;
        RECT  21.76 1.22 22.76 1.54 ;
        RECT  20.38 1.22 21.38 1.54 ;
        RECT  20.28 4.22 21.38 4.54 ;
        POLYGON  19.74 2.60 19.42 2.60 19.42 3.24 18.76 3.90 17.66 3.90
                 17.66 4.54 13.86 4.54 13.86 4.05 13.71 3.90 12.54 3.90
                 12.54 3.06 11.80 3.06 11.80 2.74 12.86 2.74 12.86 3.58
                 13.85 3.58 14.18 3.91 14.18 4.22 17.34 4.22 17.34 3.58
                 18.62 3.58 19.10 3.10 19.10 2.50 18.78 2.18 16.06 2.18
                 16.06 1.86 18.92 1.86 19.34 2.28 19.74 2.28 ;
        RECT  18.30 1.22 19.30 1.54 ;
        RECT  18.20 4.22 19.20 4.54 ;
        POLYGON  18.78 2.96 17.02 2.96 17.02 3.90 14.50 3.90 14.50 2.18
                 11.48 2.18 11.48 3.26 11.16 3.26 11.16 1.86 14.82 1.86
                 14.82 3.58 16.70 3.58 16.70 2.64 18.78 2.64 ;
        POLYGON  17.92 1.54 15.74 1.54 15.74 2.54 16.28 2.54 16.28 2.86
                 15.42 2.86 15.42 1.22 17.92 1.22 ;
        POLYGON  13.54 4.54 9.88 4.54 9.88 3.90 6.86 3.90 6.86 2.68 7.22 2.32
                 7.22 1.87 7.54 1.87 7.54 2.46 7.18 2.82 7.18 3.58 10.20 3.58
                 10.20 4.22 13.54 4.22 ;
        RECT  12.34 1.22 13.34 1.54 ;
        RECT  11.22 3.58 12.22 3.90 ;
        RECT  10.96 1.22 11.96 1.54 ;
        POLYGON  10.84 3.90 10.52 3.90 10.52 3.26 7.52 3.26 7.52 2.94
                 10.52 2.94 10.52 2.40 10.26 2.40 10.26 1.22 10.58 1.22
                 10.58 2.08 10.84 2.08 ;
        RECT  5.84 1.22 9.88 1.54 ;
        RECT  5.48 4.22 9.56 4.54 ;
        RECT  2.94 1.87 6.86 2.19 ;
        RECT  4.10 3.58 6.50 3.90 ;
        RECT  4.34 1.23 5.34 1.55 ;
        RECT  2.70 4.22 5.10 4.54 ;
        POLYGON  4.26 2.97 3.78 2.97 3.78 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 1.23 0.50 1.23 0.50 3.58 3.46 3.58 3.46 2.65 4.26 2.65 ;
        POLYGON  3.96 1.55 2.58 1.55 2.58 2.19 2.26 2.19 2.26 1.23 3.96 1.23 ;
    END
END sdffprq_4

MACRO sdffprq_2
    CLASS CORE ;
    FOREIGN sdffprq_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 26.24 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  13.52 2.72 14.18 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.65 5.28 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  25.44 3.04 25.08 3.04 25.08 4.54 24.76 4.54 24.76 1.22
                 25.08 1.22 25.08 2.72 25.44 2.72 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.44  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  8.48 2.08 8.94 2.62 ;
        END
    END rb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.60 2.65 6.34 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.65 3.04 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  26.24 0.90 25.78 0.90 25.78 1.54 25.46 1.54 25.46 0.90
                 23.46 0.90 23.46 1.54 23.14 1.54 23.14 0.90 14.04 0.90
                 14.04 1.54 13.72 1.54 13.72 0.90 1.88 0.90 1.88 1.71 0.88 1.71
                 0.88 0.90 0.00 0.90 0.00 -0.90 26.24 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  26.24 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 21.76 4.86 21.76 4.22 22.08 4.22 22.08 4.86
                 23.26 4.86 23.26 4.22 23.58 4.22 23.58 4.86 25.46 4.86
                 25.46 3.58 25.78 3.58 25.78 4.86 26.24 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  24.40 4.54 24.08 4.54 24.08 3.16 21.80 3.16 21.80 2.84
                 24.08 2.84 24.08 1.54 23.84 1.54 23.84 1.22 24.40 1.22 ;
        POLYGON  23.64 2.52 21.48 2.52 21.48 3.48 22.76 3.48 22.76 4.54
                 22.44 4.54 22.44 3.80 20.14 3.80 19.90 4.04 19.90 4.54
                 19.58 4.54 19.58 3.90 20.00 3.48 21.16 3.48 21.16 2.52
                 20.44 2.52 19.68 1.76 19.68 1.22 20.00 1.22 20.00 1.62
                 20.58 2.20 23.64 2.20 ;
        RECT  21.76 1.22 22.76 1.54 ;
        RECT  20.38 1.22 21.38 1.54 ;
        RECT  20.28 4.22 21.38 4.54 ;
        POLYGON  19.74 2.60 19.42 2.60 19.42 3.24 18.76 3.90 17.66 3.90
                 17.66 4.54 13.86 4.54 13.86 4.05 13.71 3.90 12.54 3.90
                 12.54 3.06 11.80 3.06 11.80 2.74 12.86 2.74 12.86 3.58
                 13.85 3.58 14.18 3.91 14.18 4.22 17.34 4.22 17.34 3.58
                 18.62 3.58 19.10 3.10 19.10 2.50 18.78 2.18 16.06 2.18
                 16.06 1.86 18.92 1.86 19.34 2.28 19.74 2.28 ;
        RECT  18.30 1.22 19.30 1.54 ;
        RECT  18.20 4.22 19.20 4.54 ;
        POLYGON  18.78 2.96 17.02 2.96 17.02 3.90 14.50 3.90 14.50 2.18
                 11.48 2.18 11.48 3.26 11.16 3.26 11.16 1.86 14.82 1.86
                 14.82 3.58 16.70 3.58 16.70 2.64 18.78 2.64 ;
        POLYGON  17.92 1.54 15.74 1.54 15.74 2.54 16.28 2.54 16.28 2.86
                 15.42 2.86 15.42 1.22 17.92 1.22 ;
        POLYGON  13.54 4.54 9.88 4.54 9.88 3.90 6.86 3.90 6.86 2.68 7.22 2.32
                 7.22 1.87 7.54 1.87 7.54 2.46 7.18 2.82 7.18 3.58 10.20 3.58
                 10.20 4.22 13.54 4.22 ;
        RECT  12.34 1.22 13.34 1.54 ;
        RECT  11.22 3.58 12.22 3.90 ;
        RECT  10.96 1.22 11.96 1.54 ;
        POLYGON  10.84 3.90 10.52 3.90 10.52 3.26 7.52 3.26 7.52 2.94
                 10.52 2.94 10.52 2.40 10.26 2.40 10.26 1.22 10.58 1.22
                 10.58 2.08 10.84 2.08 ;
        RECT  5.84 1.22 9.88 1.54 ;
        RECT  5.48 4.22 9.56 4.54 ;
        RECT  2.94 1.87 6.86 2.19 ;
        RECT  4.10 3.58 6.50 3.90 ;
        RECT  4.34 1.23 5.34 1.55 ;
        RECT  2.70 4.22 5.10 4.54 ;
        POLYGON  4.26 2.97 3.78 2.97 3.78 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 1.23 0.50 1.23 0.50 3.58 3.46 3.58 3.46 2.65 4.26 2.65 ;
        POLYGON  3.96 1.55 2.58 1.55 2.58 2.19 2.26 2.19 2.26 1.23 3.96 1.23 ;
    END
END sdffprq_2

MACRO sdffprq_1
    CLASS CORE ;
    FOREIGN sdffprq_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 26.24 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  13.52 2.72 14.18 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.65 5.28 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  25.44 3.04 25.08 3.04 25.08 4.54 24.76 4.54 24.76 1.22
                 25.08 1.22 25.08 2.72 25.44 2.72 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.44  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  8.48 2.08 8.94 2.62 ;
        END
    END rb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.60 2.65 6.34 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.65 3.04 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  26.24 0.90 25.78 0.90 25.78 1.54 25.46 1.54 25.46 0.90
                 23.46 0.90 23.46 1.54 23.14 1.54 23.14 0.90 14.04 0.90
                 14.04 1.14 13.72 1.14 13.72 0.90 1.88 0.90 1.88 1.71 0.88 1.71
                 0.88 0.90 0.00 0.90 0.00 -0.90 26.24 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  26.24 6.66 0.00 6.66 0.00 4.86 21.76 4.86 21.76 4.12
                 22.08 4.12 22.08 4.86 23.26 4.86 23.26 4.56 23.58 4.56
                 23.58 4.86 25.46 4.86 25.46 4.22 25.78 4.22 25.78 4.86
                 26.24 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  24.40 4.08 24.08 4.08 24.08 3.16 21.80 3.16 21.80 2.84
                 24.08 2.84 24.08 1.54 23.84 1.54 23.84 1.22 24.40 1.22 ;
        POLYGON  23.64 2.52 21.48 2.52 21.48 3.48 22.76 3.48 22.76 4.54
                 22.44 4.54 22.44 3.80 20.14 3.80 19.90 4.04 19.90 4.54
                 19.58 4.54 19.58 3.90 20.00 3.48 21.16 3.48 21.16 2.52
                 20.44 2.52 19.68 1.76 19.68 1.22 20.00 1.22 20.00 1.62
                 20.58 2.20 23.64 2.20 ;
        RECT  21.76 1.22 22.76 1.54 ;
        RECT  20.38 1.22 21.38 1.54 ;
        RECT  20.28 4.12 21.38 4.44 ;
        POLYGON  19.74 2.60 19.42 2.60 19.42 3.24 18.76 3.90 17.66 3.90
                 17.66 4.54 13.86 4.54 13.86 4.05 13.71 3.90 12.54 3.90
                 12.54 3.06 11.80 3.06 11.80 2.74 12.86 2.74 12.86 3.58
                 13.85 3.58 14.18 3.91 14.18 4.22 17.34 4.22 17.34 3.58
                 18.62 3.58 19.10 3.10 19.10 2.50 18.78 2.18 16.06 2.18
                 16.06 1.86 18.92 1.86 19.34 2.28 19.74 2.28 ;
        RECT  18.30 1.22 19.30 1.54 ;
        RECT  18.20 4.22 19.20 4.54 ;
        POLYGON  18.78 2.96 17.02 2.96 17.02 3.90 14.50 3.90 14.50 2.18
                 11.48 2.18 11.48 3.26 11.16 3.26 11.16 1.86 14.82 1.86
                 14.82 3.58 16.70 3.58 16.70 2.64 18.78 2.64 ;
        POLYGON  17.92 1.54 15.74 1.54 15.74 2.54 16.28 2.54 16.28 2.86
                 15.42 2.86 15.42 1.22 17.92 1.22 ;
        POLYGON  13.54 4.54 9.88 4.54 9.88 3.90 6.86 3.90 6.86 2.68 7.22 2.32
                 7.22 1.87 7.54 1.87 7.54 2.46 7.18 2.82 7.18 3.58 10.20 3.58
                 10.20 4.22 13.54 4.22 ;
        RECT  12.34 1.22 13.34 1.54 ;
        RECT  11.22 3.58 12.22 3.90 ;
        RECT  10.96 1.22 11.96 1.54 ;
        POLYGON  10.84 3.90 10.52 3.90 10.52 3.26 7.52 3.26 7.52 2.94
                 10.52 2.94 10.52 2.40 10.26 2.40 10.26 1.22 10.58 1.22
                 10.58 2.08 10.84 2.08 ;
        RECT  5.84 1.22 9.88 1.54 ;
        RECT  5.48 4.22 9.56 4.54 ;
        RECT  2.94 1.87 6.86 2.19 ;
        RECT  4.10 3.58 6.50 3.90 ;
        RECT  4.34 1.23 5.34 1.55 ;
        RECT  2.70 4.22 5.10 4.54 ;
        POLYGON  4.26 2.97 3.78 2.97 3.78 3.90 0.18 3.90 0.18 1.87 0.50 1.87
                 0.50 3.58 3.46 3.58 3.46 2.65 4.26 2.65 ;
        RECT  2.26 1.23 3.96 1.55 ;
    END
END sdffprq_1

MACRO sdffpr_4
    CLASS CORE ;
    FOREIGN sdffpr_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 29.44 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.86  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  29.28 3.04 28.73 3.04 28.73 4.54 26.85 4.54 26.85 4.22
                 28.41 4.22 28.41 1.54 26.85 1.54 26.85 1.22 28.73 1.22
                 28.73 2.72 29.28 2.72 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.44  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  8.48 2.08 8.94 2.62 ;
        END
    END rb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.60 2.65 6.34 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.65 3.04 3.04 ;
        END
    END se
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.35  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  26.49 3.26 24.72 3.26 24.72 1.22 26.48 1.22 26.48 1.54
                 25.04 1.54 25.04 2.72 25.44 2.72 25.44 2.94 26.49 2.94 ;
        END
    END q
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  13.52 2.72 14.18 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.65 5.28 3.04 ;
        END
    END d
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  29.44 6.66 0.00 6.66 0.00 4.86 21.76 4.86 21.76 4.12
                 22.08 4.12 22.08 4.86 23.26 4.86 23.26 4.56 23.58 4.56
                 23.58 4.86 25.46 4.86 25.46 4.52 25.78 4.52 25.78 4.86
                 29.44 4.86 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  29.44 0.90 23.46 0.90 23.46 1.54 23.14 1.54 23.14 0.90
                 14.04 0.90 14.04 1.14 13.72 1.14 13.72 0.90 1.88 0.90
                 1.88 1.71 0.88 1.71 0.88 0.90 0.00 0.90 0.00 -0.90 29.44 -0.90 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        POLYGON  28.09 2.46 27.13 2.46 27.13 3.90 24.40 3.90 24.40 4.08
                 24.08 4.08 24.08 3.16 21.80 3.16 21.80 2.84 24.08 2.84
                 24.08 1.54 23.84 1.54 23.84 1.22 24.40 1.22 24.40 3.58
                 26.81 3.58 26.81 2.14 28.09 2.14 ;
        POLYGON  23.64 2.52 21.48 2.52 21.48 3.48 22.76 3.48 22.76 4.54
                 22.44 4.54 22.44 3.80 20.14 3.80 19.90 4.04 19.90 4.54
                 19.58 4.54 19.58 3.90 20.00 3.48 21.16 3.48 21.16 2.52
                 20.44 2.52 19.68 1.76 19.68 1.22 20.00 1.22 20.00 1.62
                 20.58 2.20 23.64 2.20 ;
        RECT  21.76 1.22 22.76 1.54 ;
        RECT  20.38 1.22 21.38 1.54 ;
        RECT  20.28 4.12 21.38 4.44 ;
        POLYGON  19.74 2.60 19.42 2.60 19.42 3.24 18.76 3.90 17.66 3.90
                 17.66 4.54 13.86 4.54 13.86 4.05 13.71 3.90 12.54 3.90
                 12.54 3.06 11.80 3.06 11.80 2.74 12.86 2.74 12.86 3.58
                 13.85 3.58 14.18 3.91 14.18 4.22 17.34 4.22 17.34 3.58
                 18.62 3.58 19.10 3.10 19.10 2.50 18.78 2.18 16.06 2.18
                 16.06 1.86 18.92 1.86 19.34 2.28 19.74 2.28 ;
        RECT  18.30 1.22 19.30 1.54 ;
        RECT  18.20 4.22 19.20 4.54 ;
        POLYGON  18.78 2.96 17.02 2.96 17.02 3.90 14.50 3.90 14.50 2.18
                 11.48 2.18 11.48 3.26 11.16 3.26 11.16 1.86 14.82 1.86
                 14.82 3.58 16.70 3.58 16.70 2.64 18.78 2.64 ;
        POLYGON  17.92 1.54 15.74 1.54 15.74 2.54 16.28 2.54 16.28 2.86
                 15.42 2.86 15.42 1.22 17.92 1.22 ;
        POLYGON  13.54 4.54 9.88 4.54 9.88 3.90 6.86 3.90 6.86 2.68 7.22 2.32
                 7.22 1.87 7.54 1.87 7.54 2.46 7.18 2.82 7.18 3.58 10.20 3.58
                 10.20 4.22 13.54 4.22 ;
        RECT  12.34 1.22 13.34 1.54 ;
        RECT  11.22 3.58 12.22 3.90 ;
        RECT  10.96 1.22 11.96 1.54 ;
        POLYGON  10.84 3.90 10.52 3.90 10.52 3.26 7.52 3.26 7.52 2.94
                 10.52 2.94 10.52 2.40 10.26 2.40 10.26 1.22 10.58 1.22
                 10.58 2.08 10.84 2.08 ;
        RECT  5.84 1.22 9.88 1.54 ;
        RECT  5.48 4.22 9.56 4.54 ;
        RECT  2.94 1.87 6.86 2.19 ;
        RECT  4.10 3.58 6.50 3.90 ;
        RECT  4.34 1.23 5.34 1.55 ;
        RECT  2.70 4.22 5.10 4.54 ;
        POLYGON  4.26 2.97 3.78 2.97 3.78 3.90 0.18 3.90 0.18 1.87 0.50 1.87
                 0.50 3.58 3.46 3.58 3.46 2.65 4.26 2.65 ;
        RECT  2.26 1.23 3.96 1.55 ;
    END
END sdffpr_4

MACRO sdffpr_2
    CLASS CORE ;
    FOREIGN sdffpr_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 26.88 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  13.52 2.72 14.18 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.65 5.28 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  25.44 1.76 25.04 1.76 25.04 3.12 25.08 3.12 25.08 3.44
                 24.72 3.44 24.72 1.22 25.08 1.22 25.08 1.44 25.44 1.44 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.69  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  26.72 3.44 26.16 3.44 26.16 3.12 26.40 3.12 26.40 1.54
                 26.16 1.54 26.16 1.22 26.72 1.22 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.44  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  8.48 2.08 8.94 2.62 ;
        END
    END rb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.60 2.65 6.34 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.65 3.04 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  26.88 0.90 23.46 0.90 23.46 1.54 23.14 1.54 23.14 0.90
                 14.04 0.90 14.04 1.14 13.72 1.14 13.72 0.90 1.88 0.90
                 1.88 1.71 0.88 1.71 0.88 0.90 0.00 0.90 0.00 -0.90 26.88 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  26.88 6.66 0.00 6.66 0.00 4.86 21.76 4.86 21.76 4.12
                 22.08 4.12 22.08 4.86 23.26 4.86 23.26 4.56 23.58 4.56
                 23.58 4.86 26.88 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  25.94 2.46 25.72 2.46 25.72 4.08 24.08 4.08 24.08 3.16
                 21.80 3.16 21.80 2.84 24.08 2.84 24.08 1.54 23.84 1.54
                 23.84 1.22 24.40 1.22 24.40 3.76 25.40 3.76 25.40 2.14
                 25.94 2.14 ;
        POLYGON  23.64 2.52 21.48 2.52 21.48 3.48 22.76 3.48 22.76 4.54
                 22.44 4.54 22.44 3.80 20.14 3.80 19.90 4.04 19.90 4.54
                 19.58 4.54 19.58 3.90 20.00 3.48 21.16 3.48 21.16 2.52
                 20.44 2.52 19.68 1.76 19.68 1.22 20.00 1.22 20.00 1.62
                 20.58 2.20 23.64 2.20 ;
        RECT  21.76 1.22 22.76 1.54 ;
        RECT  20.38 1.22 21.38 1.54 ;
        RECT  20.28 4.12 21.38 4.44 ;
        POLYGON  19.74 2.60 19.42 2.60 19.42 3.24 18.76 3.90 17.66 3.90
                 17.66 4.54 13.86 4.54 13.86 4.05 13.71 3.90 12.54 3.90
                 12.54 3.06 11.80 3.06 11.80 2.74 12.86 2.74 12.86 3.58
                 13.85 3.58 14.18 3.91 14.18 4.22 17.34 4.22 17.34 3.58
                 18.62 3.58 19.10 3.10 19.10 2.50 18.78 2.18 16.06 2.18
                 16.06 1.86 18.92 1.86 19.34 2.28 19.74 2.28 ;
        RECT  18.30 1.22 19.30 1.54 ;
        RECT  18.20 4.22 19.20 4.54 ;
        POLYGON  18.78 2.96 17.02 2.96 17.02 3.90 14.50 3.90 14.50 2.18
                 11.48 2.18 11.48 3.26 11.16 3.26 11.16 1.86 14.82 1.86
                 14.82 3.58 16.70 3.58 16.70 2.64 18.78 2.64 ;
        POLYGON  17.92 1.54 15.74 1.54 15.74 2.54 16.28 2.54 16.28 2.86
                 15.42 2.86 15.42 1.22 17.92 1.22 ;
        POLYGON  13.54 4.54 9.88 4.54 9.88 3.90 6.86 3.90 6.86 2.68 7.22 2.32
                 7.22 1.87 7.54 1.87 7.54 2.46 7.18 2.82 7.18 3.58 10.20 3.58
                 10.20 4.22 13.54 4.22 ;
        RECT  12.34 1.22 13.34 1.54 ;
        RECT  11.22 3.58 12.22 3.90 ;
        RECT  10.96 1.22 11.96 1.54 ;
        POLYGON  10.84 3.90 10.52 3.90 10.52 3.26 7.52 3.26 7.52 2.94
                 10.52 2.94 10.52 2.40 10.26 2.40 10.26 1.22 10.58 1.22
                 10.58 2.08 10.84 2.08 ;
        RECT  5.84 1.22 9.88 1.54 ;
        RECT  5.48 4.22 9.56 4.54 ;
        RECT  2.94 1.87 6.86 2.19 ;
        RECT  4.10 3.58 6.50 3.90 ;
        RECT  4.34 1.23 5.34 1.55 ;
        RECT  2.70 4.22 5.10 4.54 ;
        POLYGON  4.26 2.97 3.78 2.97 3.78 3.90 0.18 3.90 0.18 1.87 0.50 1.87
                 0.50 3.58 3.46 3.58 3.46 2.65 4.26 2.65 ;
        RECT  2.26 1.23 3.96 1.55 ;
    END
END sdffpr_2

MACRO sdffpr_1
    CLASS CORE ;
    FOREIGN sdffpr_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 26.88 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  13.52 2.72 14.18 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.65 5.28 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.54  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  25.44 1.76 25.08 1.76 25.08 3.44 24.68 3.44 24.68 3.12
                 24.76 3.12 24.76 1.22 25.08 1.22 25.08 1.44 25.44 1.44 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  26.72 4.06 26.19 4.06 26.19 3.74 26.40 3.74 26.40 1.54
                 26.20 1.54 26.20 1.22 26.72 1.22 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.44  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  8.48 2.08 8.94 2.62 ;
        END
    END rb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.60 2.65 6.34 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.65 3.04 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  26.88 0.90 23.46 0.90 23.46 1.54 23.14 1.54 23.14 0.90
                 14.04 0.90 14.04 1.14 13.72 1.14 13.72 0.90 1.88 0.90
                 1.88 1.71 0.88 1.71 0.88 0.90 0.00 0.90 0.00 -0.90 26.88 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  26.88 6.66 0.00 6.66 0.00 4.86 21.76 4.86 21.76 4.12
                 22.08 4.12 22.08 4.86 23.26 4.86 23.26 4.56 23.58 4.56
                 23.58 4.86 25.50 4.86 25.50 4.56 25.82 4.56 25.82 4.86
                 26.88 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  25.98 2.46 25.72 2.46 25.72 4.08 24.04 4.08 24.04 3.16
                 21.80 3.16 21.80 2.84 24.04 2.84 24.04 1.54 23.84 1.54
                 23.84 1.22 24.36 1.22 24.36 3.76 25.40 3.76 25.40 2.14
                 25.98 2.14 ;
        POLYGON  23.64 2.52 21.48 2.52 21.48 3.48 22.76 3.48 22.76 4.54
                 22.44 4.54 22.44 3.80 20.14 3.80 19.90 4.04 19.90 4.54
                 19.58 4.54 19.58 3.90 20.00 3.48 21.16 3.48 21.16 2.52
                 20.44 2.52 19.68 1.76 19.68 1.22 20.00 1.22 20.00 1.62
                 20.58 2.20 23.64 2.20 ;
        RECT  21.76 1.22 22.76 1.54 ;
        RECT  20.38 1.22 21.38 1.54 ;
        RECT  20.28 4.12 21.38 4.44 ;
        POLYGON  19.74 2.60 19.42 2.60 19.42 3.24 18.76 3.90 17.66 3.90
                 17.66 4.54 13.86 4.54 13.86 4.05 13.71 3.90 12.54 3.90
                 12.54 3.06 11.80 3.06 11.80 2.74 12.86 2.74 12.86 3.58
                 13.85 3.58 14.18 3.91 14.18 4.22 17.34 4.22 17.34 3.58
                 18.62 3.58 19.10 3.10 19.10 2.50 18.78 2.18 16.06 2.18
                 16.06 1.86 18.92 1.86 19.34 2.28 19.74 2.28 ;
        RECT  18.30 1.22 19.30 1.54 ;
        RECT  18.20 4.22 19.20 4.54 ;
        POLYGON  18.78 2.96 17.02 2.96 17.02 3.90 14.50 3.90 14.50 2.18
                 11.48 2.18 11.48 3.26 11.16 3.26 11.16 1.86 14.82 1.86
                 14.82 3.58 16.70 3.58 16.70 2.64 18.78 2.64 ;
        POLYGON  17.92 1.54 15.74 1.54 15.74 2.54 16.28 2.54 16.28 2.86
                 15.42 2.86 15.42 1.22 17.92 1.22 ;
        POLYGON  13.54 4.54 9.88 4.54 9.88 3.90 6.86 3.90 6.86 2.68 7.22 2.32
                 7.22 1.87 7.54 1.87 7.54 2.46 7.18 2.82 7.18 3.58 10.20 3.58
                 10.20 4.22 13.54 4.22 ;
        RECT  12.34 1.22 13.34 1.54 ;
        RECT  11.22 3.58 12.22 3.90 ;
        RECT  10.96 1.22 11.96 1.54 ;
        POLYGON  10.84 3.90 10.52 3.90 10.52 3.26 7.52 3.26 7.52 2.94
                 10.52 2.94 10.52 2.40 10.26 2.40 10.26 1.22 10.58 1.22
                 10.58 2.08 10.84 2.08 ;
        RECT  5.84 1.22 9.88 1.54 ;
        RECT  5.48 4.22 9.56 4.54 ;
        RECT  2.94 1.87 6.86 2.19 ;
        RECT  4.10 3.58 6.50 3.90 ;
        RECT  4.34 1.23 5.34 1.55 ;
        RECT  2.70 4.22 5.10 4.54 ;
        POLYGON  4.26 2.97 3.78 2.97 3.78 3.90 0.18 3.90 0.18 1.87 0.50 1.87
                 0.50 3.58 3.46 3.58 3.46 2.65 4.26 2.65 ;
        RECT  2.26 1.23 3.96 1.55 ;
    END
END sdffpr_1

MACRO sdffpqb_4
    CLASS CORE ;
    FOREIGN sdffpqb_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  13.63 3.46 13.32 3.46 13.28 3.50 13.28 3.90 12.96 3.90
                 12.96 3.36 13.18 3.14 13.63 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.68 2.66 4.32 3.04 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.96 4.54 19.09 4.54 19.09 4.22 20.64 4.22 20.64 1.91
                 19.09 1.91 19.09 1.59 20.96 1.59 ;
        END
    END qb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.66 5.28 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.66 1.76 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 0.90 20.11 0.90 20.11 1.24 19.79 1.24 19.79 0.90
                 17.73 0.90 17.73 1.24 17.41 1.24 17.41 0.90 10.40 0.90
                 10.40 1.54 10.08 1.54 10.08 0.90 2.58 0.90 2.58 1.54 2.26 1.54
                 2.26 0.90 1.20 0.90 1.20 1.86 0.88 1.86 0.88 0.90 0.00 0.90
                 0.00 -0.90 21.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 10.54 4.86 10.54 3.74 10.86 3.74 10.86 4.86
                 17.53 4.86 17.53 3.96 17.85 3.96 17.85 4.86 21.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.11 3.76 18.17 3.76 18.17 3.18 17.19 3.18 17.19 2.86
                 18.17 2.86 18.17 1.22 18.49 1.22 18.49 3.44 19.79 3.44
                 19.79 2.31 20.11 2.31 ;
        POLYGON  17.85 2.47 17.53 2.47 17.53 2.28 15.63 2.28 15.63 4.54
                 15.31 4.54 15.31 2.28 14.87 1.84 14.87 1.22 15.19 1.22
                 15.19 1.70 15.45 1.96 17.85 1.96 ;
        RECT  16.09 3.96 17.09 4.28 ;
        RECT  15.69 1.22 16.99 1.54 ;
        POLYGON  14.99 3.90 13.93 3.90 13.93 3.58 14.67 3.58 14.67 2.56
                 14.29 2.18 12.11 2.18 11.89 2.40 11.89 2.58 11.57 2.58
                 11.57 2.26 11.97 1.86 14.43 1.86 14.99 2.42 ;
        RECT  11.97 4.22 14.93 4.54 ;
        RECT  11.73 1.22 14.37 1.54 ;
        POLYGON  14.13 2.82 13.04 2.82 12.44 3.42 11.69 3.42 11.69 3.90
                 11.37 3.90 11.37 3.42 10.78 3.42 10.78 2.32 8.48 2.32
                 8.48 2.00 10.78 2.00 10.78 1.22 11.10 1.22 11.10 3.10
                 12.30 3.10 12.90 2.50 14.13 2.50 ;
        RECT  9.01 3.46 10.05 3.78 ;
        RECT  8.60 1.22 9.70 1.54 ;
        POLYGON  9.69 4.54 8.30 4.54 7.66 3.90 5.72 3.90 5.72 1.86 6.04 1.86
                 6.04 3.58 7.80 3.58 8.44 4.22 9.69 4.22 ;
        POLYGON  8.63 3.63 8.31 3.63 8.31 3.26 6.38 3.26 6.38 2.94 7.80 2.94
                 7.80 1.72 7.90 1.62 7.90 1.22 8.22 1.22 8.22 1.76 8.12 1.86
                 8.12 2.94 8.63 2.94 ;
        RECT  4.34 1.22 7.52 1.54 ;
        RECT  4.34 4.22 7.52 4.54 ;
        POLYGON  5.36 2.18 1.56 2.18 1.56 1.22 1.88 1.22 1.88 1.86 5.36 1.86 ;
        RECT  2.96 3.58 5.36 3.90 ;
        RECT  2.96 1.22 3.96 1.54 ;
        RECT  1.56 4.22 3.96 4.54 ;
        POLYGON  2.74 2.98 2.40 2.98 2.40 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 1.22 0.50 1.22 0.50 3.58 2.08 3.58 2.08 2.66 2.74 2.66 ;
    END
END sdffpqb_4

MACRO sdffpqb_2
    CLASS CORE ;
    FOREIGN sdffpqb_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 20.48 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  13.63 3.46 13.32 3.46 13.28 3.50 13.28 3.90 12.96 3.90
                 12.96 3.36 13.18 3.14 13.63 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.68 2.66 4.32 3.04 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.32 4.54 19.88 4.54 19.88 4.22 20.00 4.22 20.00 1.73
                 19.55 1.73 19.55 1.41 20.32 1.41 ;
        END
    END qb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.66 5.28 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.66 1.76 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 0.90 19.17 0.90 19.17 1.24 18.85 1.24 18.85 0.90
                 17.79 0.90 17.79 1.14 17.47 1.14 17.47 0.90 10.40 0.90
                 10.40 1.54 10.08 1.54 10.08 0.90 2.58 0.90 2.58 1.54 2.26 1.54
                 2.26 0.90 1.20 0.90 1.20 1.86 0.88 1.86 0.88 0.90 0.00 0.90
                 0.00 -0.90 20.48 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 10.54 4.86 10.54 3.74 10.86 3.74 10.86 4.86
                 17.53 4.86 17.53 3.96 17.85 3.96 17.85 4.86 20.48 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  19.62 3.31 19.48 3.31 19.48 4.54 18.17 4.54 18.17 3.18
                 17.19 3.18 17.19 2.86 18.17 2.86 18.17 1.22 18.49 1.22
                 18.49 4.22 19.16 4.22 19.16 2.99 19.30 2.99 19.30 2.14
                 19.62 2.14 ;
        POLYGON  17.85 2.47 17.53 2.47 17.53 2.28 15.63 2.28 15.63 4.54
                 15.31 4.54 15.31 2.28 14.87 1.84 14.87 1.22 15.19 1.22
                 15.19 1.70 15.45 1.96 17.85 1.96 ;
        RECT  16.09 3.96 17.09 4.28 ;
        RECT  15.69 1.22 16.99 1.54 ;
        POLYGON  14.99 3.90 13.93 3.90 13.93 3.58 14.67 3.58 14.67 2.56
                 14.29 2.18 12.11 2.18 11.89 2.40 11.89 2.58 11.57 2.58
                 11.57 2.26 11.97 1.86 14.43 1.86 14.99 2.42 ;
        RECT  11.97 4.22 14.93 4.54 ;
        RECT  11.73 1.22 14.37 1.54 ;
        POLYGON  14.13 2.82 13.04 2.82 12.44 3.42 11.69 3.42 11.69 3.90
                 11.37 3.90 11.37 3.42 10.78 3.42 10.78 2.32 8.48 2.32
                 8.48 2.00 10.78 2.00 10.78 1.22 11.10 1.22 11.10 3.10
                 12.30 3.10 12.90 2.50 14.13 2.50 ;
        RECT  9.01 3.46 10.05 3.78 ;
        RECT  8.60 1.22 9.70 1.54 ;
        POLYGON  9.69 4.54 8.30 4.54 7.66 3.90 5.72 3.90 5.72 1.86 6.04 1.86
                 6.04 3.58 7.80 3.58 8.44 4.22 9.69 4.22 ;
        POLYGON  8.63 3.63 8.31 3.63 8.31 3.26 6.38 3.26 6.38 2.94 7.80 2.94
                 7.80 1.72 7.90 1.62 7.90 1.22 8.22 1.22 8.22 1.76 8.12 1.86
                 8.12 2.94 8.63 2.94 ;
        RECT  4.34 1.22 7.52 1.54 ;
        RECT  4.34 4.22 7.52 4.54 ;
        RECT  1.56 1.86 5.36 2.18 ;
        RECT  2.96 3.58 5.36 3.90 ;
        RECT  2.96 1.22 3.96 1.54 ;
        RECT  1.56 4.22 3.96 4.54 ;
        POLYGON  2.74 2.98 2.40 2.98 2.40 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 1.86 0.50 1.86 0.50 3.58 2.08 3.58 2.08 2.66 2.74 2.66 ;
    END
END sdffpqb_2

MACRO sdffpqb_1
    CLASS CORE ;
    FOREIGN sdffpqb_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 20.48 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  13.63 3.46 13.32 3.46 13.28 3.50 13.28 3.90 12.96 3.90
                 12.96 3.36 13.18 3.14 13.63 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.68 2.66 4.32 3.04 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.32 4.54 19.88 4.54 19.88 4.22 20.00 4.22 20.00 1.54
                 19.55 1.54 19.55 1.22 20.32 1.22 ;
        END
    END qb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.66 5.28 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.66 1.76 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 0.90 19.17 0.90 19.17 1.24 18.85 1.24 18.85 0.90
                 17.79 0.90 17.79 1.14 17.47 1.14 17.47 0.90 10.40 0.90
                 10.40 1.54 10.08 1.54 10.08 0.90 2.58 0.90 2.58 1.54 2.26 1.54
                 2.26 0.90 1.20 0.90 1.20 1.86 0.88 1.86 0.88 0.90 0.00 0.90
                 0.00 -0.90 20.48 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 10.54 4.86 10.54 3.74 10.86 3.74 10.86 4.86
                 17.53 4.86 17.53 3.96 17.85 3.96 17.85 4.86 20.48 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  19.62 3.95 19.48 3.95 19.48 4.54 18.17 4.54 18.17 3.18
                 17.19 3.18 17.19 2.86 18.17 2.86 18.17 1.22 18.49 1.22
                 18.49 4.22 19.16 4.22 19.16 3.63 19.30 3.63 19.30 2.14
                 19.62 2.14 ;
        POLYGON  17.85 2.47 17.53 2.47 17.53 2.28 15.63 2.28 15.63 4.54
                 15.31 4.54 15.31 2.28 14.87 1.84 14.87 1.22 15.19 1.22
                 15.19 1.70 15.45 1.96 17.85 1.96 ;
        RECT  16.09 3.96 17.09 4.28 ;
        RECT  15.69 1.22 16.99 1.54 ;
        POLYGON  14.99 3.90 13.93 3.90 13.93 3.58 14.67 3.58 14.67 2.56
                 14.29 2.18 12.11 2.18 11.89 2.40 11.89 2.58 11.57 2.58
                 11.57 2.26 11.97 1.86 14.43 1.86 14.99 2.42 ;
        RECT  11.97 4.22 14.93 4.54 ;
        RECT  11.73 1.22 14.37 1.54 ;
        POLYGON  14.13 2.82 13.04 2.82 12.44 3.42 11.69 3.42 11.69 3.90
                 11.37 3.90 11.37 3.42 10.78 3.42 10.78 2.32 8.48 2.32
                 8.48 2.00 10.78 2.00 10.78 1.22 11.10 1.22 11.10 3.10
                 12.30 3.10 12.90 2.50 14.13 2.50 ;
        RECT  9.01 3.46 10.05 3.78 ;
        RECT  8.60 1.22 9.70 1.54 ;
        POLYGON  9.69 4.54 8.30 4.54 7.66 3.90 5.72 3.90 5.72 1.86 6.04 1.86
                 6.04 3.58 7.80 3.58 8.44 4.22 9.69 4.22 ;
        POLYGON  8.63 3.63 8.31 3.63 8.31 3.26 6.38 3.26 6.38 2.94 7.80 2.94
                 7.80 1.72 7.90 1.62 7.90 1.22 8.22 1.22 8.22 1.76 8.12 1.86
                 8.12 2.94 8.63 2.94 ;
        RECT  4.34 1.22 7.52 1.54 ;
        RECT  4.34 4.22 7.52 4.54 ;
        RECT  1.56 1.86 5.36 2.18 ;
        RECT  2.96 3.58 5.36 3.90 ;
        RECT  2.96 1.22 3.96 1.54 ;
        RECT  1.56 4.22 3.96 4.54 ;
        POLYGON  2.74 2.98 2.40 2.98 2.40 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 1.86 0.50 1.86 0.50 3.58 2.08 3.58 2.08 2.66 2.74 2.66 ;
    END
END sdffpqb_1

MACRO sdffpq_4
    CLASS CORE ;
    FOREIGN sdffpq_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  13.63 3.46 13.32 3.46 13.28 3.50 13.28 3.90 12.96 3.90
                 12.96 3.36 13.18 3.14 13.63 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.68 2.66 4.32 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.76 4.54 20.44 4.54 20.44 3.04 19.36 3.04 19.36 4.54
                 19.04 4.54 19.04 3.04 18.85 3.04 18.85 1.22 19.17 1.22
                 19.17 2.72 20.25 2.72 20.25 1.22 20.57 1.22 20.57 2.72
                 20.76 2.72 ;
        END
    END q
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.66 5.28 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.66 1.76 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 0.90 19.87 0.90 19.87 1.54 19.55 1.54 19.55 0.90
                 17.74 0.90 17.74 1.14 17.42 1.14 17.42 0.90 10.40 0.90
                 10.40 1.54 10.08 1.54 10.08 0.90 2.58 0.90 2.58 1.54 2.26 1.54
                 2.26 0.90 1.20 0.90 1.20 1.40 0.88 1.40 0.88 0.90 0.00 0.90
                 0.00 -0.90 21.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 6.66 0.00 6.66 0.00 4.86 10.54 4.86 10.54 3.74
                 10.86 3.74 10.86 4.86 17.47 4.86 17.47 3.96 17.79 3.96
                 17.79 4.86 19.74 4.86 19.74 3.58 20.06 3.58 20.06 4.86
                 21.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  18.68 4.54 18.17 4.54 18.17 3.18 17.19 3.18 17.19 2.86
                 18.17 2.86 18.17 1.22 18.49 1.22 18.49 4.22 18.68 4.22 ;
        POLYGON  17.85 2.47 17.53 2.47 17.53 2.28 15.63 2.28 15.63 4.54
                 15.31 4.54 15.31 2.28 14.87 1.84 14.87 1.22 15.19 1.22
                 15.19 1.70 15.45 1.96 17.85 1.96 ;
        RECT  16.09 3.96 17.09 4.28 ;
        RECT  15.69 1.22 16.99 1.54 ;
        POLYGON  14.99 3.90 13.93 3.90 13.93 3.58 14.67 3.58 14.67 2.56
                 14.29 2.18 12.11 2.18 11.89 2.40 11.89 2.58 11.57 2.58
                 11.57 2.26 11.97 1.86 14.43 1.86 14.99 2.42 ;
        RECT  11.97 4.22 14.93 4.54 ;
        RECT  11.73 1.22 14.37 1.54 ;
        POLYGON  14.13 2.82 13.04 2.82 12.44 3.42 11.69 3.42 11.69 3.90
                 11.37 3.90 11.37 3.42 10.78 3.42 10.78 2.32 8.48 2.32
                 8.48 2.00 10.78 2.00 10.78 1.22 11.10 1.22 11.10 3.10
                 12.30 3.10 12.90 2.50 14.13 2.50 ;
        RECT  9.01 3.46 10.05 3.78 ;
        RECT  8.60 1.22 9.70 1.54 ;
        POLYGON  9.69 4.54 8.30 4.54 7.66 3.90 5.72 3.90 5.72 1.86 6.04 1.86
                 6.04 3.58 7.80 3.58 8.44 4.22 9.69 4.22 ;
        POLYGON  8.63 3.63 8.31 3.63 8.31 3.26 6.38 3.26 6.38 2.94 7.80 2.94
                 7.80 1.72 7.90 1.62 7.90 1.22 8.22 1.22 8.22 1.76 8.12 1.86
                 8.12 2.94 8.63 2.94 ;
        RECT  4.34 1.22 7.52 1.54 ;
        RECT  4.34 4.22 7.52 4.54 ;
        RECT  1.56 1.86 5.36 2.18 ;
        RECT  2.96 3.58 5.36 3.90 ;
        RECT  2.96 1.22 3.96 1.54 ;
        RECT  1.56 4.22 3.96 4.54 ;
        POLYGON  2.74 2.98 2.40 2.98 2.40 3.90 0.18 3.90 0.18 1.86 0.50 1.86
                 0.50 3.58 2.08 3.58 2.08 2.66 2.74 2.66 ;
    END
END sdffpq_4

MACRO sdffpq_2
    CLASS CORE ;
    FOREIGN sdffpq_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 20.48 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  13.63 3.46 13.32 3.46 13.28 3.50 13.28 3.90 12.96 3.90
                 12.96 3.36 13.18 3.14 13.63 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.68 2.66 4.32 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  19.68 3.04 19.36 3.04 19.36 4.54 19.04 4.54 19.04 3.04
                 18.85 3.04 18.85 1.31 19.17 1.31 19.17 2.72 19.68 2.72 ;
        END
    END q
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.66 5.28 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.66 1.76 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 0.90 19.87 0.90 19.87 1.44 19.55 1.44 19.55 0.90
                 17.74 0.90 17.74 1.14 17.42 1.14 17.42 0.90 10.40 0.90
                 10.40 1.54 10.08 1.54 10.08 0.90 2.58 0.90 2.58 1.54 2.26 1.54
                 2.26 0.90 1.20 0.90 1.20 1.40 0.88 1.40 0.88 0.90 0.00 0.90
                 0.00 -0.90 20.48 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 6.66 0.00 6.66 0.00 4.86 10.54 4.86 10.54 3.74
                 10.86 3.74 10.86 4.86 17.47 4.86 17.47 3.96 17.79 3.96
                 17.79 4.86 19.74 4.86 19.74 4.22 20.06 4.22 20.06 4.86
                 20.48 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  18.68 4.54 18.17 4.54 18.17 3.18 17.19 3.18 17.19 2.86
                 18.17 2.86 18.17 1.22 18.49 1.22 18.49 4.22 18.68 4.22 ;
        POLYGON  17.85 2.47 17.53 2.47 17.53 2.28 15.63 2.28 15.63 4.54
                 15.31 4.54 15.31 2.28 14.87 1.84 14.87 1.22 15.19 1.22
                 15.19 1.70 15.45 1.96 17.85 1.96 ;
        RECT  16.09 3.96 17.09 4.28 ;
        RECT  15.69 1.22 16.99 1.54 ;
        POLYGON  14.99 3.90 13.93 3.90 13.93 3.58 14.67 3.58 14.67 2.56
                 14.29 2.18 12.11 2.18 11.89 2.40 11.89 2.58 11.57 2.58
                 11.57 2.26 11.97 1.86 14.43 1.86 14.99 2.42 ;
        RECT  11.97 4.22 14.93 4.54 ;
        RECT  11.73 1.22 14.37 1.54 ;
        POLYGON  14.13 2.82 13.04 2.82 12.44 3.42 11.69 3.42 11.69 3.90
                 11.37 3.90 11.37 3.42 10.78 3.42 10.78 2.32 8.48 2.32
                 8.48 2.00 10.78 2.00 10.78 1.22 11.10 1.22 11.10 3.10
                 12.30 3.10 12.90 2.50 14.13 2.50 ;
        RECT  9.01 3.46 10.05 3.78 ;
        RECT  8.60 1.22 9.70 1.54 ;
        POLYGON  9.69 4.54 8.30 4.54 7.66 3.90 5.72 3.90 5.72 1.86 6.04 1.86
                 6.04 3.58 7.80 3.58 8.44 4.22 9.69 4.22 ;
        POLYGON  8.63 3.63 8.31 3.63 8.31 3.26 6.38 3.26 6.38 2.94 7.80 2.94
                 7.80 1.72 7.90 1.62 7.90 1.22 8.22 1.22 8.22 1.76 8.12 1.86
                 8.12 2.94 8.63 2.94 ;
        RECT  4.34 1.22 7.52 1.54 ;
        RECT  4.34 4.22 7.52 4.54 ;
        RECT  1.56 1.86 5.36 2.18 ;
        RECT  2.96 3.58 5.36 3.90 ;
        RECT  2.96 1.22 3.96 1.54 ;
        RECT  1.56 4.22 3.96 4.54 ;
        POLYGON  2.74 2.98 2.40 2.98 2.40 3.90 0.18 3.90 0.18 1.86 0.50 1.86
                 0.50 3.58 2.08 3.58 2.08 2.66 2.74 2.66 ;
    END
END sdffpq_2

MACRO sdffpq_1
    CLASS CORE ;
    FOREIGN sdffpq_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 20.48 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  13.63 3.46 13.32 3.46 13.28 3.50 13.28 3.90 12.96 3.90
                 12.96 3.36 13.18 3.14 13.63 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.68 2.66 4.32 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  19.68 3.04 19.36 3.04 19.36 4.30 19.04 4.30 19.04 3.04
                 18.85 3.04 18.85 1.22 19.17 1.22 19.17 2.72 19.68 2.72 ;
        END
    END q
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.66 5.28 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.66 1.76 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 0.90 19.87 0.90 19.87 1.54 19.55 1.54 19.55 0.90
                 17.74 0.90 17.74 1.14 17.42 1.14 17.42 0.90 10.40 0.90
                 10.40 1.54 10.08 1.54 10.08 0.90 2.58 0.90 2.58 1.54 2.26 1.54
                 2.26 0.90 1.20 0.90 1.20 1.86 0.88 1.86 0.88 0.90 0.00 0.90
                 0.00 -0.90 20.48 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 10.54 4.86 10.54 3.74 10.86 3.74 10.86 4.86
                 17.53 4.86 17.53 3.96 17.85 3.96 17.85 4.86 19.74 4.86
                 19.74 3.98 20.06 3.98 20.06 4.86 20.48 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  18.68 4.54 18.17 4.54 18.17 3.18 17.19 3.18 17.19 2.86
                 18.17 2.86 18.17 1.22 18.49 1.22 18.49 4.22 18.68 4.22 ;
        POLYGON  17.85 2.47 17.53 2.47 17.53 2.28 15.63 2.28 15.63 4.54
                 15.31 4.54 15.31 2.28 14.87 1.84 14.87 1.22 15.19 1.22
                 15.19 1.70 15.45 1.96 17.85 1.96 ;
        RECT  16.09 3.96 17.09 4.28 ;
        RECT  15.69 1.22 16.99 1.54 ;
        POLYGON  14.99 3.90 13.93 3.90 13.93 3.58 14.67 3.58 14.67 2.56
                 14.29 2.18 12.11 2.18 11.89 2.40 11.89 2.58 11.57 2.58
                 11.57 2.26 11.97 1.86 14.43 1.86 14.99 2.42 ;
        RECT  11.97 4.22 14.93 4.54 ;
        RECT  11.73 1.22 14.37 1.54 ;
        POLYGON  14.13 2.82 13.04 2.82 12.44 3.42 11.69 3.42 11.69 3.90
                 11.37 3.90 11.37 3.42 10.78 3.42 10.78 2.32 8.48 2.32
                 8.48 2.00 10.78 2.00 10.78 1.22 11.10 1.22 11.10 3.10
                 12.30 3.10 12.90 2.50 14.13 2.50 ;
        RECT  9.01 3.46 10.05 3.78 ;
        RECT  8.60 1.22 9.70 1.54 ;
        POLYGON  9.69 4.54 8.30 4.54 7.66 3.90 5.72 3.90 5.72 1.86 6.04 1.86
                 6.04 3.58 7.80 3.58 8.44 4.22 9.69 4.22 ;
        POLYGON  8.63 3.63 8.31 3.63 8.31 3.26 6.38 3.26 6.38 2.94 7.80 2.94
                 7.80 1.72 7.90 1.62 7.90 1.22 8.22 1.22 8.22 1.76 8.12 1.86
                 8.12 2.94 8.63 2.94 ;
        RECT  4.34 1.22 7.52 1.54 ;
        RECT  4.34 4.22 7.52 4.54 ;
        POLYGON  5.36 2.18 1.56 2.18 1.56 1.22 1.88 1.22 1.88 1.86 5.36 1.86 ;
        RECT  2.96 3.58 5.36 3.90 ;
        RECT  2.96 1.22 3.96 1.54 ;
        RECT  1.56 4.22 3.96 4.54 ;
        POLYGON  2.74 2.98 2.40 2.98 2.40 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 1.86 0.50 1.86 0.50 3.58 2.08 3.58 2.08 2.66 2.74 2.66 ;
    END
END sdffpq_1

MACRO sdffp_4
    CLASS CORE ;
    FOREIGN sdffp_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  13.63 3.46 13.32 3.46 13.28 3.50 13.28 3.90 12.96 3.90
                 12.96 3.36 13.18 3.14 13.63 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.68 2.66 4.32 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  21.10 3.26 19.33 3.26 19.33 2.94 20.64 2.94 20.64 2.72
                 20.78 2.72 20.78 1.97 18.85 1.97 18.85 1.65 21.10 1.65 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  23.52 4.54 21.42 4.54 21.42 4.22 23.20 4.22 23.20 1.91
                 21.42 1.91 21.42 1.59 23.52 1.59 ;
        END
    END qb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.66 5.28 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.66 1.76 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  23.68 0.90 22.44 0.90 22.44 1.24 22.12 1.24 22.12 0.90
                 19.87 0.90 19.87 1.25 19.55 1.25 19.55 0.90 17.73 0.90
                 17.73 1.24 17.41 1.24 17.41 0.90 10.40 0.90 10.40 1.54
                 10.08 1.54 10.08 0.90 2.58 0.90 2.58 1.54 2.26 1.54 2.26 0.90
                 1.20 0.90 1.20 1.86 0.88 1.86 0.88 0.90 0.00 0.90 0.00 -0.90
                 23.68 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  23.68 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 10.54 4.86 10.54 3.74 10.86 3.74 10.86 4.86
                 17.53 4.86 17.53 3.96 17.85 3.96 17.85 4.86 20.01 4.86
                 20.01 4.82 20.38 4.82 20.38 4.86 23.68 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  22.44 3.90 20.18 3.90 20.18 4.35 18.17 4.35 18.17 3.18
                 17.19 3.18 17.19 2.86 18.17 2.86 18.17 1.22 18.49 1.22
                 18.49 4.03 19.86 4.03 19.86 3.58 22.12 3.58 22.12 2.31
                 22.44 2.31 ;
        POLYGON  17.85 2.47 17.53 2.47 17.53 2.28 15.63 2.28 15.63 4.54
                 15.31 4.54 15.31 2.28 14.87 1.84 14.87 1.22 15.19 1.22
                 15.19 1.70 15.45 1.96 17.85 1.96 ;
        RECT  16.09 3.96 17.09 4.28 ;
        RECT  15.69 1.22 16.99 1.54 ;
        POLYGON  14.99 3.90 13.93 3.90 13.93 3.58 14.67 3.58 14.67 2.56
                 14.29 2.18 12.11 2.18 11.89 2.40 11.89 2.58 11.57 2.58
                 11.57 2.26 11.97 1.86 14.43 1.86 14.99 2.42 ;
        RECT  11.97 4.22 14.93 4.54 ;
        RECT  11.73 1.22 14.37 1.54 ;
        POLYGON  14.13 2.82 13.04 2.82 12.44 3.42 11.69 3.42 11.69 3.90
                 11.37 3.90 11.37 3.42 10.78 3.42 10.78 2.32 8.48 2.32
                 8.48 2.00 10.78 2.00 10.78 1.22 11.10 1.22 11.10 3.10
                 12.30 3.10 12.90 2.50 14.13 2.50 ;
        RECT  9.01 3.46 10.05 3.78 ;
        RECT  8.60 1.22 9.70 1.54 ;
        POLYGON  9.69 4.54 8.30 4.54 7.66 3.90 5.72 3.90 5.72 1.86 6.04 1.86
                 6.04 3.58 7.80 3.58 8.44 4.22 9.69 4.22 ;
        POLYGON  8.63 3.63 8.31 3.63 8.31 3.26 6.38 3.26 6.38 2.94 7.80 2.94
                 7.80 1.72 7.90 1.62 7.90 1.22 8.22 1.22 8.22 1.76 8.12 1.86
                 8.12 2.94 8.63 2.94 ;
        RECT  4.34 1.22 7.52 1.54 ;
        RECT  4.34 4.22 7.52 4.54 ;
        POLYGON  5.36 2.18 1.56 2.18 1.56 1.22 1.88 1.22 1.88 1.86 5.36 1.86 ;
        RECT  2.96 3.58 5.36 3.90 ;
        RECT  2.96 1.22 3.96 1.54 ;
        RECT  1.56 4.22 3.96 4.54 ;
        POLYGON  2.74 2.98 2.40 2.98 2.40 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 1.22 0.50 1.22 0.50 3.58 2.08 3.58 2.08 2.66 2.74 2.66 ;
    END
END sdffp_4

MACRO sdffp_2
    CLASS CORE ;
    FOREIGN sdffp_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  13.63 3.46 13.32 3.46 13.28 3.50 13.28 3.90 12.96 3.90
                 12.96 3.36 13.18 3.14 13.63 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.68 2.66 4.32 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.86  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  19.68 3.04 19.41 3.04 19.41 3.75 19.09 3.75 19.09 3.04
                 18.85 3.04 18.85 1.24 19.17 1.24 19.17 2.72 19.68 2.72 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.96 4.54 20.58 4.54 20.58 4.22 20.64 4.22 20.64 1.56
                 20.25 1.56 20.25 1.24 20.96 1.24 ;
        END
    END qb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.66 5.28 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.66 1.76 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 0.90 19.87 0.90 19.87 1.24 19.55 1.24 19.55 0.90
                 17.75 0.90 17.75 1.24 17.43 1.24 17.43 0.90 10.40 0.90
                 10.40 1.54 10.08 1.54 10.08 0.90 2.58 0.90 2.58 1.54 2.26 1.54
                 2.26 0.90 1.20 0.90 1.20 1.86 0.88 1.86 0.88 0.90 0.00 0.90
                 0.00 -0.90 21.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 10.54 4.86 10.54 3.74 10.86 3.74 10.86 4.86
                 17.53 4.86 17.53 3.96 17.85 3.96 17.85 4.86 21.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.32 4.00 20.18 4.00 20.18 4.54 18.17 4.54 18.17 3.18
                 17.19 3.18 17.19 2.86 18.17 2.86 18.17 1.22 18.49 1.22
                 18.49 4.22 19.86 4.22 19.86 3.68 20.00 3.68 20.00 2.14
                 20.32 2.14 ;
        POLYGON  17.85 2.47 17.53 2.47 17.53 2.28 15.63 2.28 15.63 4.54
                 15.31 4.54 15.31 2.28 14.87 1.84 14.87 1.22 15.19 1.22
                 15.19 1.70 15.45 1.96 17.85 1.96 ;
        RECT  16.09 3.96 17.09 4.28 ;
        RECT  15.69 1.22 16.99 1.54 ;
        POLYGON  14.99 3.90 13.93 3.90 13.93 3.58 14.67 3.58 14.67 2.56
                 14.29 2.18 12.11 2.18 11.89 2.40 11.89 2.58 11.57 2.58
                 11.57 2.26 11.97 1.86 14.43 1.86 14.99 2.42 ;
        RECT  11.97 4.22 14.93 4.54 ;
        RECT  11.73 1.22 14.37 1.54 ;
        POLYGON  14.13 2.82 13.04 2.82 12.44 3.42 11.69 3.42 11.69 3.90
                 11.37 3.90 11.37 3.42 10.78 3.42 10.78 2.32 8.48 2.32
                 8.48 2.00 10.78 2.00 10.78 1.22 11.10 1.22 11.10 3.10
                 12.30 3.10 12.90 2.50 14.13 2.50 ;
        RECT  9.01 3.46 10.05 3.78 ;
        RECT  8.60 1.22 9.70 1.54 ;
        POLYGON  9.69 4.54 8.30 4.54 7.66 3.90 5.72 3.90 5.72 1.86 6.04 1.86
                 6.04 3.58 7.80 3.58 8.44 4.22 9.69 4.22 ;
        POLYGON  8.63 3.63 8.31 3.63 8.31 3.26 6.38 3.26 6.38 2.94 7.80 2.94
                 7.80 1.72 7.90 1.62 7.90 1.22 8.22 1.22 8.22 1.76 8.12 1.86
                 8.12 2.94 8.63 2.94 ;
        RECT  4.34 1.22 7.52 1.54 ;
        RECT  4.34 4.22 7.52 4.54 ;
        POLYGON  5.36 2.18 1.56 2.18 1.56 1.22 1.88 1.22 1.88 1.86 5.36 1.86 ;
        RECT  2.96 3.58 5.36 3.90 ;
        RECT  2.96 1.22 3.96 1.54 ;
        RECT  1.56 4.22 3.96 4.54 ;
        POLYGON  2.74 2.98 2.40 2.98 2.40 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 1.86 0.50 1.86 0.50 3.58 2.08 3.58 2.08 2.66 2.74 2.66 ;
    END
END sdffp_2

MACRO sdffp_1
    CLASS CORE ;
    FOREIGN sdffp_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  13.63 3.46 13.32 3.46 13.28 3.50 13.28 3.90 12.96 3.90
                 12.96 3.36 13.18 3.14 13.63 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.68 2.66 4.32 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.40  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  19.68 3.04 19.41 3.04 19.41 3.90 19.09 3.90 19.09 3.04
                 18.85 3.04 18.85 1.22 19.17 1.22 19.17 2.72 19.68 2.72 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.96 4.54 20.58 4.54 20.58 4.22 20.64 4.22 20.64 1.54
                 20.25 1.54 20.25 1.22 20.96 1.22 ;
        END
    END qb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.66 5.28 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.66 1.76 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 0.90 19.87 0.90 19.87 1.24 19.55 1.24 19.55 0.90
                 17.79 0.90 17.79 1.14 17.47 1.14 17.47 0.90 10.40 0.90
                 10.40 1.54 10.08 1.54 10.08 0.90 2.58 0.90 2.58 1.54 2.26 1.54
                 2.26 0.90 1.20 0.90 1.20 1.86 0.88 1.86 0.88 0.90 0.00 0.90
                 0.00 -0.90 21.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 10.54 4.86 10.54 3.74 10.86 3.74 10.86 4.86
                 17.53 4.86 17.53 3.96 17.85 3.96 17.85 4.86 21.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.32 3.95 20.18 3.95 20.18 4.54 18.17 4.54 18.17 3.18
                 17.19 3.18 17.19 2.86 18.17 2.86 18.17 1.22 18.49 1.22
                 18.49 4.22 19.86 4.22 19.86 3.63 20.00 3.63 20.00 2.14
                 20.32 2.14 ;
        POLYGON  17.85 2.47 17.53 2.47 17.53 2.28 15.63 2.28 15.63 4.54
                 15.31 4.54 15.31 2.28 14.87 1.84 14.87 1.22 15.19 1.22
                 15.19 1.70 15.45 1.96 17.85 1.96 ;
        RECT  16.09 3.96 17.09 4.28 ;
        RECT  15.69 1.22 16.99 1.54 ;
        POLYGON  14.99 3.90 13.93 3.90 13.93 3.58 14.67 3.58 14.67 2.56
                 14.29 2.18 12.11 2.18 11.89 2.40 11.89 2.58 11.57 2.58
                 11.57 2.26 11.97 1.86 14.43 1.86 14.99 2.42 ;
        RECT  11.97 4.22 14.93 4.54 ;
        RECT  11.73 1.22 14.37 1.54 ;
        POLYGON  14.13 2.82 13.04 2.82 12.44 3.42 11.69 3.42 11.69 3.90
                 11.37 3.90 11.37 3.42 10.78 3.42 10.78 2.32 8.48 2.32
                 8.48 2.00 10.78 2.00 10.78 1.22 11.10 1.22 11.10 3.10
                 12.30 3.10 12.90 2.50 14.13 2.50 ;
        RECT  9.01 3.46 10.05 3.78 ;
        RECT  8.60 1.22 9.70 1.54 ;
        POLYGON  9.69 4.54 8.30 4.54 7.66 3.90 5.72 3.90 5.72 1.86 6.04 1.86
                 6.04 3.58 7.80 3.58 8.44 4.22 9.69 4.22 ;
        POLYGON  8.63 3.63 8.31 3.63 8.31 3.26 6.38 3.26 6.38 2.94 7.80 2.94
                 7.80 1.72 7.90 1.62 7.90 1.22 8.22 1.22 8.22 1.76 8.12 1.86
                 8.12 2.94 8.63 2.94 ;
        RECT  4.34 1.22 7.52 1.54 ;
        RECT  4.34 4.22 7.52 4.54 ;
        RECT  1.56 1.86 5.36 2.18 ;
        RECT  2.96 3.58 5.36 3.90 ;
        RECT  2.96 1.22 3.96 1.54 ;
        RECT  1.56 4.22 3.96 4.54 ;
        POLYGON  2.74 2.98 2.40 2.98 2.40 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 1.86 0.50 1.86 0.50 3.58 2.08 3.58 2.08 2.66 2.74 2.66 ;
    END
END sdffp_1

MACRO sdffnsqb_4
    CLASS CORE ;
    FOREIGN sdffnsqb_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.04 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  12.32 4.00 12.90 4.35 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.62 4.32 3.04 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  22.88 3.04 22.84 3.04 22.84 4.54 21.12 4.54 21.12 4.22
                 22.52 4.22 22.52 2.72 22.56 2.72 22.56 1.84 21.12 1.84
                 21.12 1.52 22.88 1.52 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.02  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.92 2.52 8.06 2.52 8.06 2.20 8.48 2.20 8.48 2.08 8.92 2.08 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.80 1.12 2.44 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  23.04 0.90 22.14 0.90 22.14 1.20 21.82 1.20 21.82 0.90
                 18.68 0.90 18.68 1.54 18.36 1.54 18.36 0.90 12.18 0.90
                 12.18 1.48 11.86 1.48 11.86 0.90 1.31 0.90 1.31 1.12 0.99 1.12
                 0.99 0.90 0.00 0.90 0.00 -0.90 23.04 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  23.04 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.22 1.32 4.22
                 1.32 4.86 11.44 4.86 11.44 4.16 11.76 4.16 11.76 4.86
                 14.02 4.86 14.02 4.64 14.34 4.64 14.34 4.86 17.66 4.86
                 17.66 4.62 17.98 4.62 17.98 4.86 19.74 4.86 19.74 4.00
                 20.06 4.00 20.06 4.86 23.04 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  22.14 2.48 21.40 2.48 21.40 3.12 20.76 3.12 20.76 4.54
                 20.44 4.54 20.44 3.12 19.36 3.12 19.36 4.54 19.04 4.54
                 19.04 3.12 18.18 3.12 18.18 2.80 20.44 2.80 20.44 1.52
                 20.76 1.52 20.76 2.80 21.08 2.80 21.08 2.16 22.14 2.16 ;
        POLYGON  20.12 2.48 17.86 2.48 17.86 3.64 16.50 3.64 16.50 4.48
                 16.18 4.48 16.18 3.32 17.54 3.32 17.54 2.48 16.18 2.48
                 16.18 1.22 16.50 1.22 16.50 2.16 20.12 2.16 ;
        RECT  19.06 1.22 20.06 1.54 ;
        POLYGON  18.68 4.54 18.36 4.54 18.36 4.28 17.20 4.28 17.20 4.48
                 16.88 4.48 16.88 3.96 18.36 3.96 18.36 3.58 18.68 3.58 ;
        RECT  16.88 1.22 17.98 1.54 ;
        POLYGON  15.86 3.68 11.38 3.68 11.38 3.08 9.96 3.08 9.96 2.69
                 10.28 2.69 10.28 2.76 11.70 2.76 11.70 3.36 15.54 3.36
                 15.54 2.18 14.80 2.18 14.80 1.86 15.86 1.86 ;
        POLYGON  15.80 1.54 13.56 1.54 13.56 2.18 13.24 2.18 13.24 1.22
                 15.80 1.22 ;
        RECT  13.24 4.00 15.80 4.32 ;
        POLYGON  14.56 2.92 14.36 2.92 14.36 3.04 12.35 3.04 12.35 2.44
                 10.48 2.44 10.48 2.12 12.36 2.12 12.36 1.80 12.56 1.80
                 12.56 1.24 12.88 1.24 12.88 2.12 12.68 2.12 12.68 2.72
                 14.04 2.72 14.04 2.58 14.56 2.58 ;
        RECT  10.48 1.24 11.48 1.56 ;
        RECT  10.02 3.47 11.06 3.79 ;
        POLYGON  10.70 4.54 8.68 4.54 8.68 3.90 5.96 3.90 5.96 1.86 6.28 1.86
                 6.28 3.58 9.00 3.58 9.00 4.22 10.70 4.22 ;
        POLYGON  10.10 2.18 9.64 2.18 9.64 3.90 9.32 3.90 9.32 3.16 6.60 3.16
                 6.60 2.70 6.92 2.70 6.92 2.84 9.32 2.84 9.32 1.86 9.78 1.86
                 9.78 1.22 10.10 1.22 ;
        RECT  4.58 1.22 9.40 1.54 ;
        RECT  4.58 4.22 8.36 4.54 ;
        RECT  6.66 1.86 7.66 2.18 ;
        POLYGON  5.60 2.18 1.82 2.18 1.82 1.22 2.14 1.22 2.14 1.86 5.60 1.86 ;
        RECT  2.50 3.58 5.60 3.90 ;
        RECT  2.50 1.22 4.20 1.54 ;
        RECT  1.82 4.22 4.20 4.54 ;
        POLYGON  3.00 3.08 0.48 3.08 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.76 2.68 2.76
                 2.68 2.62 3.00 2.62 ;
    END
END sdffnsqb_4

MACRO sdffnsqb_2
    CLASS CORE ;
    FOREIGN sdffnsqb_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  12.32 4.00 12.90 4.35 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.62 4.32 3.04 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  22.24 4.54 21.82 4.54 21.82 4.22 21.92 4.22 21.92 1.96
                 21.82 1.96 21.82 1.64 22.24 1.64 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.02  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.92 2.52 8.06 2.52 8.06 2.20 8.48 2.20 8.48 2.08 8.92 2.08 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.80 1.12 2.44 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  22.40 0.90 21.44 0.90 21.44 1.20 21.12 1.20 21.12 0.90
                 18.68 0.90 18.68 1.54 18.36 1.54 18.36 0.90 12.18 0.90
                 12.18 1.48 11.86 1.48 11.86 0.90 1.29 0.90 1.29 1.12 0.97 1.12
                 0.97 0.90 0.00 0.90 0.00 -0.90 22.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  22.40 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.22 1.32 4.22
                 1.32 4.86 11.44 4.86 11.44 4.16 11.76 4.16 11.76 4.86
                 14.02 4.86 14.02 4.64 14.34 4.64 14.34 4.86 17.66 4.86
                 17.66 4.62 17.98 4.62 17.98 4.86 19.74 4.86 19.74 4.22
                 20.06 4.22 20.06 4.86 21.12 4.86 21.12 3.59 21.44 3.59
                 21.44 4.86 22.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  21.54 3.12 20.76 3.12 20.76 4.54 20.44 4.54 20.44 3.12
                 19.36 3.12 19.36 4.54 19.04 4.54 19.04 3.12 18.18 3.12
                 18.18 2.80 20.34 2.80 20.34 2.16 20.40 2.16 20.40 1.22
                 20.76 1.22 20.76 1.54 20.72 1.54 20.72 2.48 20.66 2.48
                 20.66 2.80 21.22 2.80 21.22 2.36 21.54 2.36 ;
        RECT  19.06 1.22 20.06 1.54 ;
        POLYGON  20.02 2.48 17.86 2.48 17.86 3.64 16.50 3.64 16.50 4.48
                 16.18 4.48 16.18 3.32 17.54 3.32 17.54 2.48 16.18 2.48
                 16.18 1.22 16.50 1.22 16.50 2.16 20.02 2.16 ;
        POLYGON  18.68 4.54 18.36 4.54 18.36 4.28 17.20 4.28 17.20 4.48
                 16.88 4.48 16.88 3.96 18.36 3.96 18.36 3.58 18.68 3.58 ;
        RECT  16.88 1.22 17.98 1.54 ;
        POLYGON  15.86 3.68 11.38 3.68 11.38 3.08 9.96 3.08 9.96 2.69
                 10.28 2.69 10.28 2.76 11.70 2.76 11.70 3.36 15.54 3.36
                 15.54 2.18 14.80 2.18 14.80 1.86 15.86 1.86 ;
        POLYGON  15.80 1.54 13.56 1.54 13.56 2.18 13.24 2.18 13.24 1.22
                 15.80 1.22 ;
        RECT  13.24 4.00 15.80 4.32 ;
        POLYGON  14.56 2.92 14.36 2.92 14.36 3.04 12.35 3.04 12.35 2.44
                 10.48 2.44 10.48 2.12 12.36 2.12 12.36 1.80 12.56 1.80
                 12.56 1.58 12.88 1.58 12.88 2.12 12.68 2.12 12.68 2.72
                 14.04 2.72 14.04 2.58 14.56 2.58 ;
        RECT  10.48 1.24 11.48 1.56 ;
        RECT  10.02 3.47 11.06 3.79 ;
        POLYGON  10.70 4.54 8.68 4.54 8.68 3.90 5.96 3.90 5.96 1.86 6.28 1.86
                 6.28 3.58 9.00 3.58 9.00 4.22 10.70 4.22 ;
        POLYGON  10.10 2.18 9.64 2.18 9.64 3.90 9.32 3.90 9.32 3.16 6.60 3.16
                 6.60 2.70 6.92 2.70 6.92 2.84 9.32 2.84 9.32 1.86 9.78 1.86
                 9.78 1.22 10.10 1.22 ;
        RECT  4.58 1.22 9.40 1.54 ;
        RECT  4.58 4.22 8.36 4.54 ;
        RECT  6.66 1.86 7.66 2.18 ;
        POLYGON  5.60 2.18 1.82 2.18 1.82 1.22 2.14 1.22 2.14 1.86 5.60 1.86 ;
        RECT  2.50 3.58 5.60 3.90 ;
        RECT  2.50 1.22 4.20 1.54 ;
        POLYGON  4.20 4.54 1.82 4.54 1.82 3.58 2.14 3.58 2.14 4.22 4.20 4.22 ;
        POLYGON  3.00 3.08 0.48 3.08 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.76 2.68 2.76
                 2.68 2.62 3.00 2.62 ;
    END
END sdffnsqb_2

MACRO sdffnsqb_1
    CLASS CORE ;
    FOREIGN sdffnsqb_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  12.32 4.00 12.90 4.35 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.62 4.32 3.04 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  22.24 4.54 21.82 4.54 21.82 4.22 21.92 4.22 21.92 1.54
                 21.82 1.54 21.82 1.22 22.24 1.22 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.02  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.92 2.52 8.06 2.52 8.06 2.20 8.48 2.20 8.48 2.08 8.92 2.08 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.80 1.12 2.44 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  22.40 0.90 21.44 0.90 21.44 1.20 21.12 1.20 21.12 0.90
                 18.68 0.90 18.68 1.54 18.36 1.54 18.36 0.90 12.18 0.90
                 12.18 1.48 11.86 1.48 11.86 0.90 1.29 0.90 1.29 1.12 0.97 1.12
                 0.97 0.90 0.00 0.90 0.00 -0.90 22.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  22.40 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.22 1.32 4.22
                 1.32 4.86 11.44 4.86 11.44 4.16 11.76 4.16 11.76 4.86
                 14.02 4.86 14.02 4.64 14.34 4.64 14.34 4.86 17.66 4.86
                 17.66 4.62 17.98 4.62 17.98 4.86 19.74 4.86 19.74 4.22
                 20.06 4.22 20.06 4.86 21.12 4.86 21.12 3.75 21.44 3.75
                 21.44 4.86 22.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  21.54 3.12 20.76 3.12 20.76 4.54 20.44 4.54 20.44 3.12
                 19.36 3.12 19.36 4.54 19.04 4.54 19.04 3.12 18.18 3.12
                 18.18 2.80 20.34 2.80 20.34 2.16 20.40 2.16 20.40 1.22
                 20.76 1.22 20.76 1.54 20.72 1.54 20.72 2.48 20.66 2.48
                 20.66 2.80 21.22 2.80 21.22 2.36 21.54 2.36 ;
        RECT  19.06 1.22 20.06 1.54 ;
        POLYGON  20.02 2.48 17.86 2.48 17.86 3.64 16.50 3.64 16.50 4.48
                 16.18 4.48 16.18 3.32 17.54 3.32 17.54 2.48 16.18 2.48
                 16.18 1.22 16.50 1.22 16.50 2.16 20.02 2.16 ;
        POLYGON  18.68 4.54 18.36 4.54 18.36 4.28 17.20 4.28 17.20 4.48
                 16.88 4.48 16.88 3.96 18.36 3.96 18.36 3.58 18.68 3.58 ;
        RECT  16.88 1.22 17.98 1.54 ;
        POLYGON  15.86 3.68 11.38 3.68 11.38 3.08 9.96 3.08 9.96 2.69
                 10.28 2.69 10.28 2.76 11.70 2.76 11.70 3.36 15.54 3.36
                 15.54 2.18 14.80 2.18 14.80 1.86 15.86 1.86 ;
        POLYGON  15.80 1.54 13.56 1.54 13.56 2.18 13.24 2.18 13.24 1.22
                 15.80 1.22 ;
        RECT  13.24 4.00 15.80 4.32 ;
        POLYGON  14.56 2.92 14.36 2.92 14.36 3.04 12.35 3.04 12.35 2.44
                 10.48 2.44 10.48 2.12 12.36 2.12 12.36 1.80 12.56 1.80
                 12.56 1.58 12.88 1.58 12.88 2.12 12.68 2.12 12.68 2.72
                 14.04 2.72 14.04 2.58 14.56 2.58 ;
        RECT  10.48 1.24 11.48 1.56 ;
        RECT  10.02 3.47 11.06 3.79 ;
        POLYGON  10.70 4.54 8.68 4.54 8.68 3.90 5.96 3.90 5.96 1.86 6.28 1.86
                 6.28 3.58 9.00 3.58 9.00 4.22 10.70 4.22 ;
        POLYGON  10.10 2.18 9.64 2.18 9.64 3.90 9.32 3.90 9.32 3.16 6.60 3.16
                 6.60 2.70 6.92 2.70 6.92 2.84 9.32 2.84 9.32 1.86 9.78 1.86
                 9.78 1.22 10.10 1.22 ;
        RECT  4.58 1.22 9.40 1.54 ;
        RECT  4.58 4.22 8.36 4.54 ;
        RECT  6.66 1.86 7.66 2.18 ;
        POLYGON  5.60 2.18 1.82 2.18 1.82 1.22 2.14 1.22 2.14 1.86 5.60 1.86 ;
        RECT  2.50 3.58 5.60 3.90 ;
        RECT  2.50 1.22 4.20 1.54 ;
        POLYGON  4.20 4.54 1.82 4.54 1.82 3.58 2.14 3.58 2.14 4.22 4.20 4.22 ;
        POLYGON  3.00 3.08 0.48 3.08 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.76 2.68 2.76
                 2.68 2.62 3.00 2.62 ;
    END
END sdffnsqb_1

MACRO sdffnsq_4
    CLASS CORE ;
    FOREIGN sdffnsq_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.04 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  12.32 4.00 12.90 4.35 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.62 4.32 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  22.84 4.54 22.52 4.54 22.52 3.04 21.44 3.04 21.44 4.54
                 21.12 4.54 21.12 1.22 21.44 1.22 21.44 2.72 22.52 2.72
                 22.52 1.22 22.84 1.22 ;
        END
    END q
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.02  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.92 2.52 8.06 2.52 8.06 2.20 8.48 2.20 8.48 2.08 8.92 2.08 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.80 1.12 2.44 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  23.04 0.90 22.14 0.90 22.14 1.54 21.82 1.54 21.82 0.90
                 18.68 0.90 18.68 1.54 18.36 1.54 18.36 0.90 12.18 0.90
                 12.18 1.48 11.86 1.48 11.86 0.90 1.31 0.90 1.31 1.12 0.99 1.12
                 0.99 0.90 0.00 0.90 0.00 -0.90 23.04 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  23.04 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.22 1.32 4.22
                 1.32 4.86 11.44 4.86 11.44 4.16 11.76 4.16 11.76 4.86
                 14.02 4.86 14.02 4.64 14.34 4.64 14.34 4.86 17.66 4.86
                 17.66 4.62 17.98 4.62 17.98 4.86 19.74 4.86 19.74 4.00
                 20.06 4.00 20.06 4.86 21.82 4.86 21.82 3.58 22.14 3.58
                 22.14 4.86 23.04 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.76 4.54 20.44 4.54 20.44 3.12 19.36 3.12 19.36 4.54
                 19.04 4.54 19.04 3.12 18.18 3.12 18.18 2.80 20.44 2.80
                 20.44 1.22 20.76 1.22 ;
        POLYGON  20.12 2.48 17.86 2.48 17.86 3.64 16.50 3.64 16.50 4.48
                 16.18 4.48 16.18 3.32 17.54 3.32 17.54 2.48 16.18 2.48
                 16.18 1.22 16.50 1.22 16.50 2.16 20.12 2.16 ;
        RECT  19.06 1.22 20.06 1.54 ;
        POLYGON  18.68 4.54 18.36 4.54 18.36 4.28 17.20 4.28 17.20 4.48
                 16.88 4.48 16.88 3.96 18.36 3.96 18.36 3.58 18.68 3.58 ;
        RECT  16.88 1.22 17.98 1.54 ;
        POLYGON  15.86 3.68 11.38 3.68 11.38 3.08 9.96 3.08 9.96 2.69
                 10.28 2.69 10.28 2.76 11.70 2.76 11.70 3.36 15.54 3.36
                 15.54 2.18 14.80 2.18 14.80 1.86 15.86 1.86 ;
        POLYGON  15.80 1.54 13.56 1.54 13.56 2.18 13.24 2.18 13.24 1.22
                 15.80 1.22 ;
        RECT  13.24 4.00 15.80 4.32 ;
        POLYGON  14.56 2.92 14.36 2.92 14.36 3.04 12.35 3.04 12.35 2.44
                 10.48 2.44 10.48 2.12 12.36 2.12 12.36 1.80 12.56 1.80
                 12.56 1.24 12.88 1.24 12.88 2.12 12.68 2.12 12.68 2.72
                 14.04 2.72 14.04 2.58 14.56 2.58 ;
        RECT  10.48 1.24 11.48 1.56 ;
        RECT  10.02 3.47 11.06 3.79 ;
        POLYGON  10.70 4.54 8.68 4.54 8.68 3.90 5.96 3.90 5.96 1.86 6.28 1.86
                 6.28 3.58 9.00 3.58 9.00 4.22 10.70 4.22 ;
        POLYGON  10.10 2.18 9.64 2.18 9.64 3.90 9.32 3.90 9.32 3.16 6.60 3.16
                 6.60 2.70 6.92 2.70 6.92 2.84 9.32 2.84 9.32 1.86 9.78 1.86
                 9.78 1.22 10.10 1.22 ;
        RECT  4.58 1.22 9.40 1.54 ;
        RECT  4.58 4.22 8.36 4.54 ;
        RECT  6.66 1.86 7.66 2.18 ;
        POLYGON  5.60 2.18 1.82 2.18 1.82 1.22 2.14 1.22 2.14 1.86 5.60 1.86 ;
        RECT  2.50 3.58 5.60 3.90 ;
        RECT  2.50 1.22 4.20 1.54 ;
        POLYGON  4.20 4.54 1.82 4.54 1.82 3.58 2.14 3.58 2.14 4.22 4.20 4.22 ;
        POLYGON  3.00 3.08 0.48 3.08 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.76 2.68 2.76
                 2.68 2.62 3.00 2.62 ;
    END
END sdffnsq_4

MACRO sdffnsq_2
    CLASS CORE ;
    FOREIGN sdffnsq_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  12.32 4.00 12.90 4.35 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.62 4.32 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  22.24 3.04 22.14 3.04 22.14 4.54 21.82 4.54 21.82 1.22
                 22.14 1.22 22.14 2.72 22.24 2.72 ;
        END
    END q
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.02  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.92 2.52 8.06 2.52 8.06 2.20 8.48 2.20 8.48 2.08 8.92 2.08 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.80 1.12 2.44 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  22.40 0.90 21.44 0.90 21.44 1.54 21.12 1.54 21.12 0.90
                 18.68 0.90 18.68 1.54 18.36 1.54 18.36 0.90 12.18 0.90
                 12.18 1.48 11.86 1.48 11.86 0.90 1.32 0.90 1.32 1.12 1.00 1.12
                 1.00 0.90 0.00 0.90 0.00 -0.90 22.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  22.40 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.22 1.32 4.22
                 1.32 4.86 11.44 4.86 11.44 4.16 11.76 4.16 11.76 4.86
                 14.02 4.86 14.02 4.64 14.34 4.64 14.34 4.86 17.66 4.86
                 17.66 4.62 17.98 4.62 17.98 4.86 19.74 4.86 19.74 4.00
                 20.06 4.00 20.06 4.86 21.12 4.86 21.12 3.58 21.44 3.58
                 21.44 4.86 22.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.76 4.54 20.44 4.54 20.44 3.12 19.36 3.12 19.36 4.54
                 19.04 4.54 19.04 3.12 18.18 3.12 18.18 2.80 20.44 2.80
                 20.44 1.22 20.76 1.22 ;
        POLYGON  20.12 2.48 17.86 2.48 17.86 3.64 16.50 3.64 16.50 4.48
                 16.18 4.48 16.18 3.32 17.54 3.32 17.54 2.48 16.18 2.48
                 16.18 1.22 16.50 1.22 16.50 2.16 20.12 2.16 ;
        RECT  19.06 1.22 20.06 1.54 ;
        POLYGON  18.68 4.54 18.36 4.54 18.36 4.28 17.20 4.28 17.20 4.48
                 16.88 4.48 16.88 3.96 18.36 3.96 18.36 3.58 18.68 3.58 ;
        RECT  16.88 1.22 17.98 1.54 ;
        POLYGON  15.86 3.68 11.38 3.68 11.38 3.08 9.96 3.08 9.96 2.69
                 10.28 2.69 10.28 2.76 11.70 2.76 11.70 3.36 15.54 3.36
                 15.54 2.18 14.80 2.18 14.80 1.86 15.86 1.86 ;
        POLYGON  15.80 1.54 13.56 1.54 13.56 2.18 13.24 2.18 13.24 1.22
                 15.80 1.22 ;
        RECT  13.24 4.00 15.80 4.32 ;
        POLYGON  14.56 2.92 14.36 2.92 14.36 3.04 12.35 3.04 12.35 2.44
                 10.48 2.44 10.48 2.12 12.36 2.12 12.36 1.80 12.56 1.80
                 12.56 1.24 12.88 1.24 12.88 2.12 12.68 2.12 12.68 2.72
                 14.04 2.72 14.04 2.58 14.56 2.58 ;
        RECT  10.48 1.24 11.48 1.56 ;
        RECT  10.02 3.47 11.06 3.79 ;
        POLYGON  10.70 4.54 8.68 4.54 8.68 3.90 5.96 3.90 5.96 1.86 6.28 1.86
                 6.28 3.58 9.00 3.58 9.00 4.22 10.70 4.22 ;
        POLYGON  10.10 2.18 9.64 2.18 9.64 3.90 9.32 3.90 9.32 3.16 6.60 3.16
                 6.60 2.70 6.92 2.70 6.92 2.84 9.32 2.84 9.32 1.86 9.78 1.86
                 9.78 1.22 10.10 1.22 ;
        RECT  4.58 1.22 9.40 1.54 ;
        RECT  4.58 4.22 8.36 4.54 ;
        RECT  6.66 1.86 7.66 2.18 ;
        POLYGON  5.60 2.18 1.82 2.18 1.82 1.22 2.14 1.22 2.14 1.86 5.60 1.86 ;
        RECT  2.50 3.58 5.60 3.90 ;
        RECT  2.50 1.22 4.20 1.54 ;
        POLYGON  4.20 4.54 1.82 4.54 1.82 3.58 2.14 3.58 2.14 4.22 4.20 4.22 ;
        POLYGON  3.00 3.08 0.48 3.08 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.76 2.68 2.76
                 2.68 2.62 3.00 2.62 ;
    END
END sdffnsq_2

MACRO sdffnsq_1
    CLASS CORE ;
    FOREIGN sdffnsq_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  12.32 4.00 12.90 4.35 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.62 4.32 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  22.24 3.04 22.14 3.04 22.14 4.54 21.82 4.54 21.82 1.22
                 22.14 1.22 22.14 2.72 22.24 2.72 ;
        END
    END q
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.02  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.92 2.52 8.06 2.52 8.06 2.20 8.48 2.20 8.48 2.08 8.92 2.08 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.80 1.12 2.44 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  22.40 0.90 21.44 0.90 21.44 1.54 21.12 1.54 21.12 0.90
                 18.68 0.90 18.68 1.54 18.36 1.54 18.36 0.90 12.18 0.90
                 12.18 1.56 11.86 1.56 11.86 0.90 1.29 0.90 1.29 1.12 0.97 1.12
                 0.97 0.90 0.00 0.90 0.00 -0.90 22.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  22.40 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.22 1.32 4.22
                 1.32 4.86 11.44 4.86 11.44 4.16 11.76 4.16 11.76 4.86
                 14.02 4.86 14.02 4.64 14.34 4.64 14.34 4.86 17.66 4.86
                 17.66 4.62 17.98 4.62 17.98 4.86 19.74 4.86 19.74 4.00
                 20.06 4.00 20.06 4.86 21.12 4.86 21.12 4.22 21.44 4.22
                 21.44 4.86 22.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.76 4.54 20.44 4.54 20.44 3.12 19.36 3.12 19.36 4.54
                 19.04 4.54 19.04 3.12 18.18 3.12 18.18 2.80 20.44 2.80
                 20.44 1.22 20.76 1.22 ;
        POLYGON  20.12 2.48 17.86 2.48 17.86 3.64 16.50 3.64 16.50 4.48
                 16.18 4.48 16.18 3.32 17.54 3.32 17.54 2.48 16.18 2.48
                 16.18 1.22 16.50 1.22 16.50 2.16 20.12 2.16 ;
        RECT  19.06 1.22 20.06 1.54 ;
        POLYGON  18.68 4.54 18.36 4.54 18.36 4.28 17.20 4.28 17.20 4.48
                 16.88 4.48 16.88 3.96 18.36 3.96 18.36 3.58 18.68 3.58 ;
        RECT  16.88 1.22 17.98 1.54 ;
        POLYGON  15.86 3.68 11.38 3.68 11.38 3.08 9.96 3.08 9.96 2.69
                 10.28 2.69 10.28 2.76 11.70 2.76 11.70 3.36 15.54 3.36
                 15.54 2.18 14.80 2.18 14.80 1.86 15.86 1.86 ;
        POLYGON  15.80 1.54 13.56 1.54 13.56 2.18 13.24 2.18 13.24 1.22
                 15.80 1.22 ;
        RECT  13.24 4.00 15.80 4.32 ;
        POLYGON  14.56 2.92 14.36 2.92 14.36 3.04 12.35 3.04 12.35 2.44
                 10.48 2.44 10.48 2.12 12.35 2.12 12.35 1.84 12.56 1.84
                 12.56 1.24 12.88 1.24 12.88 2.16 12.67 2.16 12.67 2.72
                 14.04 2.72 14.04 2.58 14.56 2.58 ;
        RECT  10.48 1.24 11.48 1.56 ;
        RECT  10.02 3.47 11.06 3.79 ;
        POLYGON  10.70 4.54 8.68 4.54 8.68 3.90 5.96 3.90 5.96 1.86 6.28 1.86
                 6.28 3.58 9.00 3.58 9.00 4.22 10.70 4.22 ;
        POLYGON  10.10 2.18 9.64 2.18 9.64 3.90 9.32 3.90 9.32 3.16 6.60 3.16
                 6.60 2.70 6.92 2.70 6.92 2.84 9.32 2.84 9.32 1.86 9.78 1.86
                 9.78 1.22 10.10 1.22 ;
        RECT  4.58 1.22 9.40 1.54 ;
        RECT  4.58 4.22 8.36 4.54 ;
        RECT  6.66 1.86 7.66 2.18 ;
        POLYGON  5.60 2.18 1.82 2.18 1.82 1.22 2.14 1.22 2.14 1.86 5.60 1.86 ;
        RECT  2.50 3.58 5.60 3.90 ;
        RECT  2.50 1.22 4.20 1.54 ;
        RECT  1.82 4.22 4.20 4.54 ;
        POLYGON  3.00 3.08 0.48 3.08 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.76 2.68 2.76
                 2.68 2.62 3.00 2.62 ;
    END
END sdffnsq_1

MACRO sdffns_4
    CLASS CORE ;
    FOREIGN sdffns_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 25.60 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  12.32 4.00 12.90 4.35 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.62 4.32 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  22.84 1.84 21.44 1.84 21.44 2.72 21.60 2.72 21.60 2.94
                 22.84 2.94 22.84 3.26 21.12 3.26 21.12 1.52 22.84 1.52 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  25.44 3.04 24.92 3.04 24.92 4.54 23.20 4.54 23.20 4.22
                 24.60 4.22 24.60 2.72 24.74 2.72 24.74 1.84 23.20 1.84
                 23.20 1.52 25.06 1.52 25.06 2.72 25.44 2.72 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.02  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.92 2.52 8.06 2.52 8.06 2.20 8.48 2.20 8.48 2.08 8.92 2.08 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.80 1.12 2.44 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  25.60 0.90 24.22 0.90 24.22 1.20 23.90 1.20 23.90 0.90
                 22.14 0.90 22.14 1.20 21.82 1.20 21.82 0.90 18.68 0.90
                 18.68 1.54 18.36 1.54 18.36 0.90 12.18 0.90 12.18 1.48
                 11.86 1.48 11.86 0.90 1.31 0.90 1.31 1.12 0.99 1.12 0.99 0.90
                 0.00 0.90 0.00 -0.90 25.60 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  25.60 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.22 1.32 4.22
                 1.32 4.86 11.44 4.86 11.44 4.16 11.76 4.16 11.76 4.86
                 14.02 4.86 14.02 4.64 14.34 4.64 14.34 4.86 17.66 4.86
                 17.66 4.62 17.98 4.62 17.98 4.86 19.74 4.86 19.74 4.00
                 20.06 4.00 20.06 4.86 21.82 4.86 21.82 4.22 22.14 4.22
                 22.14 4.86 25.60 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  24.22 2.48 23.48 2.48 23.48 3.90 20.76 3.90 20.76 4.54
                 20.44 4.54 20.44 3.12 19.36 3.12 19.36 4.54 19.04 4.54
                 19.04 3.12 18.18 3.12 18.18 2.80 20.44 2.80 20.44 1.52
                 20.76 1.52 20.76 3.58 23.16 3.58 23.16 2.16 24.22 2.16 ;
        POLYGON  20.12 2.48 17.86 2.48 17.86 3.64 16.50 3.64 16.50 4.48
                 16.18 4.48 16.18 3.32 17.54 3.32 17.54 2.48 16.18 2.48
                 16.18 1.22 16.50 1.22 16.50 2.16 20.12 2.16 ;
        RECT  19.06 1.22 20.06 1.54 ;
        POLYGON  18.68 4.54 18.36 4.54 18.36 4.28 17.20 4.28 17.20 4.48
                 16.88 4.48 16.88 3.96 18.36 3.96 18.36 3.58 18.68 3.58 ;
        RECT  16.88 1.22 17.98 1.54 ;
        POLYGON  15.86 3.68 11.38 3.68 11.38 3.08 9.96 3.08 9.96 2.69
                 10.28 2.69 10.28 2.76 11.70 2.76 11.70 3.36 15.54 3.36
                 15.54 2.18 14.80 2.18 14.80 1.86 15.86 1.86 ;
        POLYGON  15.80 1.54 13.56 1.54 13.56 2.18 13.24 2.18 13.24 1.22
                 15.80 1.22 ;
        RECT  13.24 4.00 15.80 4.32 ;
        POLYGON  14.56 2.92 14.36 2.92 14.36 3.04 12.35 3.04 12.35 2.44
                 10.48 2.44 10.48 2.12 12.36 2.12 12.36 1.80 12.56 1.80
                 12.56 1.24 12.88 1.24 12.88 2.12 12.68 2.12 12.68 2.72
                 14.04 2.72 14.04 2.58 14.56 2.58 ;
        RECT  10.48 1.24 11.48 1.56 ;
        RECT  10.02 3.47 11.06 3.79 ;
        POLYGON  10.70 4.54 8.68 4.54 8.68 3.90 5.96 3.90 5.96 1.86 6.28 1.86
                 6.28 3.58 9.00 3.58 9.00 4.22 10.70 4.22 ;
        POLYGON  10.10 2.18 9.64 2.18 9.64 3.90 9.32 3.90 9.32 3.16 6.60 3.16
                 6.60 2.70 6.92 2.70 6.92 2.84 9.32 2.84 9.32 1.86 9.78 1.86
                 9.78 1.22 10.10 1.22 ;
        RECT  4.58 1.22 9.40 1.54 ;
        RECT  4.58 4.22 8.36 4.54 ;
        RECT  6.66 1.86 7.66 2.18 ;
        POLYGON  5.60 2.18 1.82 2.18 1.82 1.22 2.14 1.22 2.14 1.86 5.60 1.86 ;
        RECT  2.50 3.58 5.60 3.90 ;
        RECT  2.50 1.22 4.20 1.54 ;
        RECT  1.82 4.22 4.20 4.54 ;
        POLYGON  3.00 3.08 0.48 3.08 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.76 2.68 2.76
                 2.68 2.62 3.00 2.62 ;
    END
END sdffns_4

MACRO sdffns_2
    CLASS CORE ;
    FOREIGN sdffns_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.04 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  12.32 4.00 12.90 4.35 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.62 4.32 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.77  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  21.60 3.04 21.44 3.04 21.44 3.26 20.98 3.26 20.98 2.94
                 21.12 2.94 21.12 1.22 21.44 1.22 21.44 2.72 21.60 2.72 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  22.88 4.54 22.52 4.54 22.52 4.22 22.56 4.22 22.56 1.54
                 22.52 1.54 22.52 1.22 22.88 1.22 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.02  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.92 2.52 8.06 2.52 8.06 2.20 8.48 2.20 8.48 2.08 8.92 2.08 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.80 1.12 2.44 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  23.04 0.90 22.14 0.90 22.14 1.54 21.82 1.54 21.82 0.90
                 18.68 0.90 18.68 1.54 18.36 1.54 18.36 0.90 12.18 0.90
                 12.18 1.48 11.86 1.48 11.86 0.90 1.29 0.90 1.29 1.12 0.97 1.12
                 0.97 0.90 0.00 0.90 0.00 -0.90 23.04 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  23.04 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.22 1.32 4.22
                 1.32 4.86 11.44 4.86 11.44 4.16 11.76 4.16 11.76 4.86
                 14.02 4.86 14.02 4.64 14.34 4.64 14.34 4.86 17.66 4.86
                 17.66 4.62 17.98 4.62 17.98 4.86 19.74 4.86 19.74 4.22
                 20.06 4.22 20.06 4.86 21.82 4.86 21.82 4.22 22.14 4.22
                 22.14 4.86 23.04 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  22.24 3.90 20.76 3.90 20.76 4.54 20.44 4.54 20.44 3.90
                 20.34 3.90 20.34 3.12 19.36 3.12 19.36 4.54 19.04 4.54
                 19.04 3.12 18.18 3.12 18.18 2.80 20.34 2.80 20.34 2.16
                 20.40 2.16 20.40 1.22 20.76 1.22 20.76 1.54 20.72 1.54
                 20.72 2.48 20.66 2.48 20.66 3.58 21.92 3.58 21.92 2.40
                 22.24 2.40 ;
        RECT  19.06 1.22 20.06 1.54 ;
        POLYGON  20.02 2.48 17.86 2.48 17.86 3.64 16.50 3.64 16.50 4.48
                 16.18 4.48 16.18 3.32 17.54 3.32 17.54 2.48 16.18 2.48
                 16.18 1.22 16.50 1.22 16.50 2.16 20.02 2.16 ;
        POLYGON  18.68 4.54 18.36 4.54 18.36 4.28 17.20 4.28 17.20 4.48
                 16.88 4.48 16.88 3.96 18.36 3.96 18.36 3.58 18.68 3.58 ;
        RECT  16.88 1.22 17.98 1.54 ;
        POLYGON  15.86 3.68 11.38 3.68 11.38 3.08 9.96 3.08 9.96 2.69
                 10.28 2.69 10.28 2.76 11.70 2.76 11.70 3.36 15.54 3.36
                 15.54 2.18 14.80 2.18 14.80 1.86 15.86 1.86 ;
        RECT  13.24 1.22 15.80 1.54 ;
        RECT  13.24 4.00 15.80 4.32 ;
        POLYGON  14.56 2.92 14.36 2.92 14.36 3.04 12.35 3.04 12.35 2.44
                 10.48 2.44 10.48 2.12 12.36 2.12 12.36 1.80 12.56 1.80
                 12.56 1.58 12.88 1.58 12.88 2.12 12.68 2.12 12.68 2.72
                 14.04 2.72 14.04 2.58 14.56 2.58 ;
        RECT  10.48 1.24 11.48 1.56 ;
        RECT  10.02 3.47 11.06 3.79 ;
        POLYGON  10.70 4.54 8.68 4.54 8.68 3.90 5.96 3.90 5.96 1.86 6.28 1.86
                 6.28 3.58 9.00 3.58 9.00 4.22 10.70 4.22 ;
        POLYGON  10.10 2.18 9.64 2.18 9.64 3.90 9.32 3.90 9.32 3.16 6.60 3.16
                 6.60 2.70 6.92 2.70 6.92 2.84 9.32 2.84 9.32 1.86 9.78 1.86
                 9.78 1.22 10.10 1.22 ;
        RECT  4.58 1.22 9.40 1.54 ;
        RECT  4.58 4.22 8.36 4.54 ;
        RECT  6.66 1.86 7.66 2.18 ;
        POLYGON  5.60 2.18 1.82 2.18 1.82 1.22 2.14 1.22 2.14 1.86 5.60 1.86 ;
        RECT  2.50 3.58 5.60 3.90 ;
        RECT  2.50 1.22 4.20 1.54 ;
        POLYGON  4.20 4.54 1.82 4.54 1.82 3.58 2.14 3.58 2.14 4.22 4.20 4.22 ;
        POLYGON  3.00 3.08 0.48 3.08 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.76 2.68 2.76
                 2.68 2.62 3.00 2.62 ;
    END
END sdffns_2

MACRO sdffns_1
    CLASS CORE ;
    FOREIGN sdffns_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.04 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  12.32 4.00 12.90 4.35 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.62 4.32 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.30  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  21.60 3.04 21.44 3.04 21.44 3.26 20.98 3.26 20.98 2.94
                 21.12 2.94 21.12 1.22 21.44 1.22 21.44 2.72 21.60 2.72 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  22.88 4.54 22.52 4.54 22.52 4.22 22.56 4.22 22.56 1.54
                 22.52 1.54 22.52 1.22 22.88 1.22 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.02  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.92 2.52 8.06 2.52 8.06 2.20 8.48 2.20 8.48 2.08 8.92 2.08 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.80 1.12 2.44 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  23.04 0.90 22.14 0.90 22.14 1.20 21.82 1.20 21.82 0.90
                 18.68 0.90 18.68 1.54 18.36 1.54 18.36 0.90 12.18 0.90
                 12.18 1.48 11.86 1.48 11.86 0.90 1.29 0.90 1.29 1.12 0.97 1.12
                 0.97 0.90 0.00 0.90 0.00 -0.90 23.04 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  23.04 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.22 1.32 4.22
                 1.32 4.86 11.44 4.86 11.44 4.16 11.76 4.16 11.76 4.86
                 14.02 4.86 14.02 4.64 14.34 4.64 14.34 4.86 17.66 4.86
                 17.66 4.62 17.98 4.62 17.98 4.86 19.74 4.86 19.74 4.22
                 20.06 4.22 20.06 4.86 21.82 4.86 21.82 4.38 22.14 4.38
                 22.14 4.86 23.04 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  22.24 3.90 20.76 3.90 20.76 4.54 20.44 4.54 20.44 3.90
                 20.34 3.90 20.34 3.12 19.36 3.12 19.36 4.54 19.04 4.54
                 19.04 3.12 18.18 3.12 18.18 2.80 20.34 2.80 20.34 2.16
                 20.40 2.16 20.40 1.22 20.76 1.22 20.76 1.54 20.72 1.54
                 20.72 2.48 20.66 2.48 20.66 3.58 21.92 3.58 21.92 2.40
                 22.24 2.40 ;
        RECT  19.06 1.22 20.06 1.54 ;
        POLYGON  20.02 2.48 17.86 2.48 17.86 3.64 16.50 3.64 16.50 4.48
                 16.18 4.48 16.18 3.32 17.54 3.32 17.54 2.48 16.18 2.48
                 16.18 1.22 16.50 1.22 16.50 2.16 20.02 2.16 ;
        POLYGON  18.68 4.54 18.36 4.54 18.36 4.28 17.20 4.28 17.20 4.48
                 16.88 4.48 16.88 3.96 18.36 3.96 18.36 3.58 18.68 3.58 ;
        RECT  16.88 1.22 17.98 1.54 ;
        POLYGON  15.86 3.68 11.38 3.68 11.38 3.08 9.96 3.08 9.96 2.69
                 10.28 2.69 10.28 2.76 11.70 2.76 11.70 3.36 15.54 3.36
                 15.54 2.18 14.80 2.18 14.80 1.86 15.86 1.86 ;
        POLYGON  15.80 1.54 13.56 1.54 13.56 2.18 13.24 2.18 13.24 1.22
                 15.80 1.22 ;
        RECT  13.24 4.00 15.80 4.32 ;
        POLYGON  14.56 2.92 14.36 2.92 14.36 3.04 12.35 3.04 12.35 2.44
                 10.48 2.44 10.48 2.12 12.36 2.12 12.36 1.80 12.56 1.80
                 12.56 1.58 12.88 1.58 12.88 2.12 12.68 2.12 12.68 2.72
                 14.04 2.72 14.04 2.58 14.56 2.58 ;
        RECT  10.48 1.24 11.48 1.56 ;
        RECT  10.02 3.47 11.06 3.79 ;
        POLYGON  10.70 4.54 8.68 4.54 8.68 3.90 5.96 3.90 5.96 1.86 6.28 1.86
                 6.28 3.58 9.00 3.58 9.00 4.22 10.70 4.22 ;
        POLYGON  10.10 2.18 9.64 2.18 9.64 3.90 9.32 3.90 9.32 3.16 6.60 3.16
                 6.60 2.70 6.92 2.70 6.92 2.84 9.32 2.84 9.32 1.86 9.78 1.86
                 9.78 1.22 10.10 1.22 ;
        RECT  4.58 1.22 9.40 1.54 ;
        RECT  4.58 4.22 8.36 4.54 ;
        RECT  6.66 1.86 7.66 2.18 ;
        POLYGON  5.60 2.18 1.82 2.18 1.82 1.22 2.14 1.22 2.14 1.86 5.60 1.86 ;
        RECT  2.50 3.58 5.60 3.90 ;
        RECT  2.50 1.22 4.20 1.54 ;
        POLYGON  4.20 4.54 1.82 4.54 1.82 3.58 2.14 3.58 2.14 4.22 4.20 4.22 ;
        POLYGON  3.00 3.08 0.48 3.08 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.76 2.68 2.76
                 2.68 2.62 3.00 2.62 ;
    END
END sdffns_1

MACRO sdffnrsqb_4
    CLASS CORE ;
    FOREIGN sdffnrsqb_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 28.16 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.96 3.04 15.84 3.04 15.84 2.72 16.64 2.72 16.64 2.50
                 16.96 2.50 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.62 4.56 3.04 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.97  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  26.91 1.54 26.84 1.54 26.84 4.47 26.52 4.47 26.52 1.76
                 26.40 1.76 26.40 1.22 26.91 1.22 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.52 3.04 6.80 3.04 6.80 2.60 7.20 2.60 7.20 2.72 7.52 2.72 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  23.16 2.62 23.52 3.24 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.95 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.76 1.12 2.40 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  28.16 0.90 25.97 0.90 25.97 1.52 25.65 1.52 25.65 0.90
                 23.01 0.90 23.01 1.53 22.69 1.53 22.69 0.90 1.33 0.90
                 1.33 1.12 1.01 1.12 1.01 0.90 0.00 0.90 0.00 -0.90 28.16 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  28.16 6.66 0.00 6.66 0.00 4.86 1.02 4.86 1.02 4.22 1.34 4.22
                 1.34 4.86 3.24 4.86 3.24 4.66 3.56 4.66 3.56 4.86 15.22 4.86
                 15.22 4.14 15.54 4.14 15.54 4.64 17.98 4.64 17.98 4.86
                 21.14 4.86 21.14 4.60 21.46 4.60 21.46 4.86 25.70 4.86
                 25.70 3.62 26.02 3.62 26.02 4.86 27.22 4.86 27.22 4.25
                 27.54 4.25 27.54 4.86 28.16 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  26.13 2.57 25.27 2.57 25.27 3.90 22.84 3.90 22.84 4.54
                 22.52 4.54 22.52 3.58 22.25 3.58 22.25 3.26 22.84 3.26
                 22.84 3.58 24.95 3.58 24.95 1.22 25.27 1.22 25.27 2.25
                 26.13 2.25 ;
        RECT  23.27 4.22 25.20 4.54 ;
        RECT  23.57 1.22 24.57 1.54 ;
        POLYGON  24.16 2.64 23.84 2.64 23.84 2.24 21.93 2.24 21.93 3.64
                 20.08 3.64 20.08 4.54 19.76 4.54 19.76 3.32 21.61 3.32
                 21.61 2.24 20.19 2.24 20.19 1.28 20.51 1.28 20.51 1.92
                 24.16 1.92 ;
        RECT  20.89 1.28 22.21 1.60 ;
        POLYGON  22.16 4.28 20.78 4.28 20.78 4.44 20.46 4.44 20.46 3.96
                 22.16 3.96 ;
        POLYGON  19.81 1.60 19.49 1.60 19.49 1.54 17.17 1.54 17.17 1.22
                 19.81 1.22 ;
        POLYGON  19.46 3.20 18.70 3.20 18.70 3.68 18.38 3.68 18.38 2.88
                 18.81 2.88 18.81 2.18 16.45 2.18 16.45 1.54 14.62 1.54
                 14.62 2.40 13.48 2.40 13.48 2.08 14.30 2.08 14.30 1.22
                 16.77 1.22 16.77 1.86 19.13 1.86 19.13 2.88 19.46 2.88 ;
        RECT  16.80 4.00 19.38 4.32 ;
        POLYGON  18.06 3.08 17.88 3.08 17.88 3.68 16.44 3.68 16.44 4.32
                 16.12 4.32 16.12 3.68 15.00 3.68 15.00 3.06 12.52 3.06
                 12.52 2.52 12.84 2.52 12.84 2.74 15.00 2.74 15.00 1.86
                 16.13 1.86 16.13 2.18 15.32 2.18 15.32 3.36 17.56 3.36
                 17.56 2.76 18.06 2.76 ;
        POLYGON  14.68 3.90 13.68 3.90 13.68 3.46 14.00 3.46 14.00 3.58
                 14.68 3.58 ;
        POLYGON  14.16 4.54 11.78 4.54 11.24 4.00 11.24 3.26 8.52 3.26
                 7.74 2.48 7.74 1.86 8.06 1.86 8.06 2.34 8.66 2.94 11.56 2.94
                 11.56 3.86 11.92 4.22 14.16 4.22 ;
        RECT  12.82 1.28 13.98 1.60 ;
        POLYGON  13.30 3.90 12.06 3.90 11.88 3.72 11.88 2.62 9.76 2.62
                 9.76 2.30 11.88 2.30 11.88 1.96 11.98 1.86 12.08 1.86
                 12.08 1.28 12.40 1.28 12.40 2.18 12.20 2.18 12.20 3.58
                 13.30 3.58 ;
        POLYGON  11.70 1.60 11.38 1.60 11.38 1.54 4.62 1.54 4.62 1.22
                 11.70 1.22 ;
        RECT  4.62 4.22 11.00 4.54 ;
        RECT  7.76 3.58 10.32 3.90 ;
        RECT  8.46 1.86 9.46 2.18 ;
        POLYGON  7.26 2.20 6.94 2.20 6.94 2.18 6.32 2.18 6.32 3.90 6.00 3.90
                 6.00 1.86 7.26 1.86 ;
        POLYGON  5.64 2.18 1.86 2.18 1.86 1.22 2.18 1.22 2.18 1.86 5.64 1.86 ;
        POLYGON  5.64 3.72 5.32 3.72 5.32 3.70 2.54 3.70 2.54 3.38 5.64 3.38 ;
        RECT  2.54 1.22 4.24 1.54 ;
        POLYGON  4.24 4.34 1.86 4.34 1.86 3.38 2.18 3.38 2.18 4.02 4.24 4.02 ;
        POLYGON  3.24 3.04 0.48 3.04 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.72 2.92 2.72
                 2.92 2.60 3.24 2.60 ;
    END
END sdffnrsqb_4

MACRO sdffnrsqb_2
    CLASS CORE ;
    FOREIGN sdffnrsqb_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 27.52 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.96 3.04 15.84 3.04 15.84 2.72 16.64 2.72 16.64 2.50
                 16.96 2.50 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.62 4.56 3.04 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.84  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  27.36 2.40 26.88 2.40 26.88 3.06 26.92 3.06 26.92 3.38
                 26.56 3.38 26.56 1.22 26.91 1.22 26.91 1.54 26.88 1.54
                 26.88 2.08 27.36 2.08 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.52 3.04 6.80 3.04 6.80 2.60 7.20 2.60 7.20 2.72 7.52 2.72 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  23.16 2.62 23.52 3.26 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.95 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.76 1.12 2.40 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  27.52 0.90 25.97 0.90 25.97 1.52 25.65 1.52 25.65 0.90
                 23.01 0.90 23.01 1.53 22.69 1.53 22.69 0.90 1.32 0.90
                 1.32 1.12 1.00 1.12 1.00 0.90 0.00 0.90 0.00 -0.90 27.52 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  27.52 6.66 0.00 6.66 0.00 4.86 1.03 4.86 1.03 4.22 1.35 4.22
                 1.35 4.86 3.24 4.86 3.24 4.66 3.56 4.66 3.56 4.86 15.22 4.86
                 15.22 4.14 15.54 4.14 15.54 4.64 17.98 4.64 17.98 4.86
                 21.14 4.86 21.14 4.60 21.46 4.60 21.46 4.86 27.52 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  26.13 2.57 25.27 2.57 25.27 3.90 22.84 3.90 22.84 4.54
                 22.52 4.54 22.52 3.58 22.25 3.58 22.25 3.26 22.84 3.26
                 22.84 3.58 24.95 3.58 24.95 1.22 25.27 1.22 25.27 2.25
                 26.13 2.25 ;
        RECT  23.27 4.22 25.20 4.54 ;
        RECT  23.57 1.22 24.57 1.54 ;
        POLYGON  24.16 2.64 23.84 2.64 23.84 2.24 21.93 2.24 21.93 3.64
                 20.08 3.64 20.08 4.54 19.76 4.54 19.76 3.32 21.61 3.32
                 21.61 2.24 20.19 2.24 20.19 1.28 20.51 1.28 20.51 1.92
                 24.16 1.92 ;
        RECT  20.89 1.28 22.21 1.60 ;
        POLYGON  22.16 4.28 20.78 4.28 20.78 4.44 20.46 4.44 20.46 3.96
                 22.16 3.96 ;
        POLYGON  19.81 1.60 19.49 1.60 19.49 1.54 17.17 1.54 17.17 1.22
                 19.81 1.22 ;
        POLYGON  19.46 3.20 18.70 3.20 18.70 3.68 18.38 3.68 18.38 2.88
                 18.81 2.88 18.81 2.18 16.45 2.18 16.45 1.54 14.62 1.54
                 14.62 2.40 13.48 2.40 13.48 2.08 14.30 2.08 14.30 1.22
                 16.77 1.22 16.77 1.86 19.13 1.86 19.13 2.88 19.46 2.88 ;
        RECT  16.80 4.00 19.38 4.32 ;
        POLYGON  18.06 3.08 17.88 3.08 17.88 3.68 16.44 3.68 16.44 4.32
                 16.12 4.32 16.12 3.68 15.00 3.68 15.00 3.06 12.52 3.06
                 12.52 2.52 12.84 2.52 12.84 2.74 15.00 2.74 15.00 1.86
                 16.13 1.86 16.13 2.18 15.32 2.18 15.32 3.36 17.56 3.36
                 17.56 2.76 18.06 2.76 ;
        POLYGON  14.68 3.90 13.68 3.90 13.68 3.46 14.00 3.46 14.00 3.58
                 14.68 3.58 ;
        POLYGON  14.16 4.54 11.78 4.54 11.24 4.00 11.24 3.26 8.52 3.26
                 7.74 2.48 7.74 1.86 8.06 1.86 8.06 2.34 8.66 2.94 11.56 2.94
                 11.56 3.86 11.92 4.22 14.16 4.22 ;
        RECT  12.82 1.28 13.98 1.60 ;
        POLYGON  13.30 3.90 12.06 3.90 11.88 3.72 11.88 2.62 9.76 2.62
                 9.76 2.30 11.88 2.30 11.88 1.96 11.98 1.86 12.08 1.86
                 12.08 1.28 12.40 1.28 12.40 2.18 12.20 2.18 12.20 3.58
                 13.30 3.58 ;
        POLYGON  11.70 1.60 11.38 1.60 11.38 1.54 4.62 1.54 4.62 1.22
                 11.70 1.22 ;
        RECT  4.62 4.22 11.00 4.54 ;
        RECT  7.76 3.58 10.32 3.90 ;
        RECT  8.46 1.86 9.46 2.18 ;
        POLYGON  7.26 2.20 6.94 2.20 6.94 2.18 6.32 2.18 6.32 3.90 6.00 3.90
                 6.00 1.86 7.26 1.86 ;
        POLYGON  5.64 2.18 1.86 2.18 1.86 1.22 2.18 1.22 2.18 1.86 5.64 1.86 ;
        POLYGON  5.64 3.72 5.32 3.72 5.32 3.70 2.54 3.70 2.54 3.38 5.64 3.38 ;
        RECT  2.54 1.22 4.24 1.54 ;
        POLYGON  4.24 4.34 1.86 4.34 1.86 3.38 2.18 3.38 2.18 4.02 4.24 4.02 ;
        POLYGON  3.24 3.04 0.48 3.04 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.72 2.92 2.72
                 2.92 2.60 3.24 2.60 ;
    END
END sdffnrsqb_2

MACRO sdffnrsqb_1
    CLASS CORE ;
    FOREIGN sdffnrsqb_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 27.52 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.96 3.04 15.84 3.04 15.84 2.72 16.64 2.72 16.64 2.50
                 16.96 2.50 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.62 4.56 3.04 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.56  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  27.36 2.40 26.88 2.40 26.88 3.06 26.92 3.06 26.92 3.38
                 26.56 3.38 26.56 1.22 26.91 1.22 26.91 1.54 26.88 1.54
                 26.88 2.08 27.36 2.08 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.52 3.04 6.80 3.04 6.80 2.60 7.20 2.60 7.20 2.72 7.52 2.72 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  23.16 2.62 23.52 3.26 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.95 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.76 1.12 2.40 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  27.52 0.90 26.10 0.90 26.10 1.52 25.78 1.52 25.78 0.90
                 23.01 0.90 23.01 1.53 22.69 1.53 22.69 0.90 1.32 0.90
                 1.32 1.12 1.00 1.12 1.00 0.90 0.00 0.90 0.00 -0.90 27.52 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  27.52 6.66 0.00 6.66 0.00 4.86 0.99 4.86 0.99 4.22 1.31 4.22
                 1.31 4.86 3.24 4.86 3.24 4.66 3.56 4.66 3.56 4.86 15.22 4.86
                 15.22 4.14 15.54 4.14 15.54 4.64 17.98 4.64 17.98 4.86
                 21.14 4.86 21.14 4.60 21.46 4.60 21.46 4.86 27.52 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  26.13 2.57 25.27 2.57 25.27 3.90 22.84 3.90 22.84 4.54
                 22.52 4.54 22.52 3.58 22.25 3.58 22.25 3.26 22.84 3.26
                 22.84 3.58 24.95 3.58 24.95 1.22 25.27 1.22 25.27 2.25
                 26.13 2.25 ;
        RECT  23.27 4.22 25.20 4.54 ;
        RECT  23.57 1.22 24.57 1.54 ;
        POLYGON  24.16 2.64 23.84 2.64 23.84 2.24 21.93 2.24 21.93 3.64
                 20.08 3.64 20.08 4.54 19.76 4.54 19.76 3.32 21.61 3.32
                 21.61 2.24 20.19 2.24 20.19 1.28 20.51 1.28 20.51 1.92
                 24.16 1.92 ;
        RECT  20.89 1.28 22.21 1.60 ;
        POLYGON  22.16 4.28 20.78 4.28 20.78 4.44 20.46 4.44 20.46 3.96
                 22.16 3.96 ;
        POLYGON  19.81 1.60 19.49 1.60 19.49 1.54 17.17 1.54 17.17 1.22
                 19.81 1.22 ;
        POLYGON  19.46 3.20 18.70 3.20 18.70 3.68 18.38 3.68 18.38 2.88
                 18.81 2.88 18.81 2.18 16.45 2.18 16.45 1.54 14.62 1.54
                 14.62 2.40 13.48 2.40 13.48 2.08 14.30 2.08 14.30 1.22
                 16.77 1.22 16.77 1.86 19.13 1.86 19.13 2.88 19.46 2.88 ;
        RECT  16.80 4.00 19.38 4.32 ;
        POLYGON  18.06 3.08 17.88 3.08 17.88 3.68 16.44 3.68 16.44 4.32
                 16.12 4.32 16.12 3.68 15.00 3.68 15.00 3.06 12.52 3.06
                 12.52 2.52 12.84 2.52 12.84 2.74 15.00 2.74 15.00 1.86
                 16.13 1.86 16.13 2.18 15.32 2.18 15.32 3.36 17.56 3.36
                 17.56 2.76 18.06 2.76 ;
        POLYGON  14.68 3.90 13.68 3.90 13.68 3.46 14.00 3.46 14.00 3.58
                 14.68 3.58 ;
        POLYGON  14.16 4.54 11.78 4.54 11.24 4.00 11.24 3.26 8.52 3.26
                 7.74 2.48 7.74 1.86 8.06 1.86 8.06 2.34 8.66 2.94 11.56 2.94
                 11.56 3.86 11.92 4.22 14.16 4.22 ;
        RECT  12.82 1.28 13.98 1.60 ;
        POLYGON  13.30 3.90 12.06 3.90 11.88 3.72 11.88 2.62 9.76 2.62
                 9.76 2.30 11.88 2.30 11.88 1.96 11.98 1.86 12.08 1.86
                 12.08 1.28 12.40 1.28 12.40 2.18 12.20 2.18 12.20 3.58
                 13.30 3.58 ;
        POLYGON  11.70 1.60 11.38 1.60 11.38 1.54 4.62 1.54 4.62 1.22
                 11.70 1.22 ;
        RECT  4.62 4.22 11.00 4.54 ;
        RECT  7.76 3.58 10.32 3.90 ;
        RECT  8.46 1.86 9.46 2.18 ;
        POLYGON  7.26 2.20 6.94 2.20 6.94 2.18 6.32 2.18 6.32 3.90 6.00 3.90
                 6.00 1.86 7.26 1.86 ;
        POLYGON  5.64 2.18 1.86 2.18 1.86 1.22 2.18 1.22 2.18 1.86 5.64 1.86 ;
        POLYGON  5.64 3.72 5.32 3.72 5.32 3.70 2.54 3.70 2.54 3.38 5.64 3.38 ;
        RECT  2.54 1.22 4.24 1.54 ;
        POLYGON  4.24 4.34 1.86 4.34 1.86 3.38 2.18 3.38 2.18 4.02 4.24 4.02 ;
        POLYGON  3.24 3.04 0.48 3.04 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.72 2.92 2.72
                 2.92 2.60 3.24 2.60 ;
    END
END sdffnrsqb_1

MACRO sdffnrsq_4
    CLASS CORE ;
    FOREIGN sdffnrsq_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 29.44 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.96 3.04 15.84 3.04 15.84 2.72 16.64 2.72 16.64 2.50
                 16.96 2.50 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.62 4.56 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  29.00 3.28 28.99 3.28 28.99 4.54 28.67 4.54 28.67 2.40
                 27.74 2.40 27.74 3.28 27.59 3.28 27.59 4.54 27.27 4.54
                 27.27 2.96 27.42 2.96 27.42 1.54 27.27 1.54 27.27 1.22
                 27.74 1.22 27.74 2.08 28.67 2.08 28.67 1.22 29.00 1.22 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.52 3.04 6.80 3.04 6.80 2.60 7.20 2.60 7.20 2.72 7.52 2.72 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  23.16 2.62 23.52 3.26 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.95 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.76 1.12 2.40 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  29.44 0.90 25.97 0.90 25.97 1.52 25.65 1.52 25.65 0.90
                 23.01 0.90 23.01 1.53 22.69 1.53 22.69 0.90 1.33 0.90
                 1.33 1.12 1.01 1.12 1.01 0.90 0.00 0.90 0.00 -0.90 29.44 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  29.44 6.66 0.00 6.66 0.00 4.86 1.02 4.86 1.02 4.22 1.34 4.22
                 1.34 4.86 3.24 4.86 3.24 4.66 3.56 4.66 3.56 4.86 15.22 4.86
                 15.22 4.14 15.54 4.14 15.54 4.64 17.98 4.64 17.98 4.86
                 21.14 4.86 21.14 4.60 21.46 4.60 21.46 4.86 25.70 4.86
                 25.70 3.58 26.02 3.58 26.02 4.86 27.97 4.86 27.97 3.58
                 28.29 3.58 28.29 4.86 29.44 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  27.07 2.46 26.88 2.46 26.88 4.54 26.56 4.54 26.56 1.22
                 26.91 1.22 26.91 1.54 26.88 1.54 26.88 2.14 27.07 2.14 ;
        POLYGON  26.13 2.57 25.27 2.57 25.27 3.90 22.84 3.90 22.84 4.54
                 22.52 4.54 22.52 3.58 22.25 3.58 22.25 3.26 22.84 3.26
                 22.84 3.58 24.95 3.58 24.95 1.22 25.27 1.22 25.27 2.25
                 26.13 2.25 ;
        RECT  23.27 4.22 25.20 4.54 ;
        RECT  23.57 1.22 24.57 1.54 ;
        POLYGON  24.16 2.64 23.84 2.64 23.84 2.24 21.93 2.24 21.93 3.64
                 20.08 3.64 20.08 4.54 19.76 4.54 19.76 3.32 21.61 3.32
                 21.61 2.24 20.19 2.24 20.19 1.28 20.51 1.28 20.51 1.92
                 24.16 1.92 ;
        RECT  20.89 1.28 22.21 1.60 ;
        POLYGON  22.16 4.28 20.78 4.28 20.78 4.44 20.46 4.44 20.46 3.96
                 22.16 3.96 ;
        POLYGON  19.81 1.60 19.49 1.60 19.49 1.54 17.17 1.54 17.17 1.22
                 19.81 1.22 ;
        POLYGON  19.46 3.20 18.70 3.20 18.70 3.68 18.38 3.68 18.38 2.88
                 18.81 2.88 18.81 2.18 16.45 2.18 16.45 1.54 14.62 1.54
                 14.62 2.40 13.48 2.40 13.48 2.08 14.30 2.08 14.30 1.22
                 16.77 1.22 16.77 1.86 19.13 1.86 19.13 2.88 19.46 2.88 ;
        RECT  16.80 4.00 19.38 4.32 ;
        POLYGON  18.06 3.08 17.88 3.08 17.88 3.68 16.44 3.68 16.44 4.32
                 16.12 4.32 16.12 3.68 15.00 3.68 15.00 3.06 12.52 3.06
                 12.52 2.52 12.84 2.52 12.84 2.74 15.00 2.74 15.00 1.86
                 16.13 1.86 16.13 2.18 15.32 2.18 15.32 3.36 17.56 3.36
                 17.56 2.76 18.06 2.76 ;
        POLYGON  14.68 3.90 13.68 3.90 13.68 3.46 14.00 3.46 14.00 3.58
                 14.68 3.58 ;
        POLYGON  14.16 4.54 11.78 4.54 11.24 4.00 11.24 3.26 8.52 3.26
                 7.74 2.48 7.74 1.86 8.06 1.86 8.06 2.34 8.66 2.94 11.56 2.94
                 11.56 3.86 11.92 4.22 14.16 4.22 ;
        RECT  12.82 1.28 13.98 1.60 ;
        POLYGON  13.30 3.90 12.06 3.90 11.88 3.72 11.88 2.62 9.76 2.62
                 9.76 2.30 11.88 2.30 11.88 1.96 11.98 1.86 12.08 1.86
                 12.08 1.28 12.40 1.28 12.40 2.18 12.20 2.18 12.20 3.58
                 13.30 3.58 ;
        POLYGON  11.70 1.60 11.38 1.60 11.38 1.54 4.62 1.54 4.62 1.22
                 11.70 1.22 ;
        RECT  4.62 4.22 11.00 4.54 ;
        RECT  7.76 3.58 10.32 3.90 ;
        RECT  8.46 1.86 9.46 2.18 ;
        POLYGON  7.26 2.20 6.94 2.20 6.94 2.18 6.32 2.18 6.32 3.90 6.00 3.90
                 6.00 1.86 7.26 1.86 ;
        POLYGON  5.64 2.18 1.86 2.18 1.86 1.22 2.18 1.22 2.18 1.86 5.64 1.86 ;
        POLYGON  5.64 3.72 5.32 3.72 5.32 3.70 2.54 3.70 2.54 3.38 5.64 3.38 ;
        RECT  2.54 1.22 4.24 1.54 ;
        POLYGON  4.24 4.34 1.86 4.34 1.86 3.38 2.18 3.38 2.18 4.02 4.24 4.02 ;
        POLYGON  3.24 3.04 0.48 3.04 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.72 2.92 2.72
                 2.92 2.60 3.24 2.60 ;
    END
END sdffnrsq_4

MACRO sdffnrsq_2
    CLASS CORE ;
    FOREIGN sdffnrsq_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 28.80 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.96 3.04 15.84 3.04 15.84 2.72 16.64 2.72 16.64 2.50
                 16.96 2.50 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.62 4.56 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  28.00 2.40 27.74 2.40 27.74 3.28 27.59 3.28 27.59 4.54
                 27.27 4.54 27.27 2.96 27.42 2.96 27.42 1.66 27.27 1.66
                 27.27 1.34 27.74 1.34 27.74 2.08 28.00 2.08 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.52 3.04 6.80 3.04 6.80 2.60 7.20 2.60 7.20 2.72 7.52 2.72 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  23.16 2.62 23.52 3.26 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.95 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.76 1.12 2.40 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  28.80 0.90 26.09 0.90 26.09 1.52 25.77 1.52 25.77 0.90
                 23.01 0.90 23.01 1.53 22.69 1.53 22.69 0.90 1.33 0.90
                 1.33 1.12 1.01 1.12 1.01 0.90 0.00 0.90 0.00 -0.90 28.80 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  28.80 6.66 0.00 6.66 0.00 4.86 1.02 4.86 1.02 4.22 1.34 4.22
                 1.34 4.86 3.24 4.86 3.24 4.66 3.56 4.66 3.56 4.86 15.22 4.86
                 15.22 4.14 15.54 4.14 15.54 4.64 17.98 4.64 17.98 4.86
                 21.14 4.86 21.14 4.60 21.46 4.60 21.46 4.86 25.70 4.86
                 25.70 4.22 26.02 4.22 26.02 4.86 27.97 4.86 27.97 3.75
                 28.29 3.75 28.29 4.86 28.80 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  27.07 2.46 26.88 2.46 26.88 4.54 26.56 4.54 26.56 1.22
                 26.91 1.22 26.91 1.54 26.88 1.54 26.88 2.14 27.07 2.14 ;
        POLYGON  26.13 2.57 25.27 2.57 25.27 3.90 22.84 3.90 22.84 4.54
                 22.52 4.54 22.52 3.58 22.25 3.58 22.25 3.26 22.84 3.26
                 22.84 3.58 24.95 3.58 24.95 1.22 25.27 1.22 25.27 2.25
                 26.13 2.25 ;
        RECT  23.27 4.22 25.20 4.54 ;
        RECT  23.57 1.22 24.57 1.54 ;
        POLYGON  24.16 2.64 23.84 2.64 23.84 2.24 21.93 2.24 21.93 3.64
                 20.08 3.64 20.08 4.54 19.76 4.54 19.76 3.32 21.61 3.32
                 21.61 2.24 20.19 2.24 20.19 1.28 20.51 1.28 20.51 1.92
                 24.16 1.92 ;
        RECT  20.89 1.28 22.21 1.60 ;
        POLYGON  22.16 4.28 20.78 4.28 20.78 4.44 20.46 4.44 20.46 3.96
                 22.16 3.96 ;
        POLYGON  19.81 1.60 19.49 1.60 19.49 1.54 17.17 1.54 17.17 1.22
                 19.81 1.22 ;
        POLYGON  19.46 3.20 18.70 3.20 18.70 3.68 18.38 3.68 18.38 2.88
                 18.81 2.88 18.81 2.18 16.45 2.18 16.45 1.54 14.62 1.54
                 14.62 2.40 13.48 2.40 13.48 2.08 14.30 2.08 14.30 1.22
                 16.77 1.22 16.77 1.86 19.13 1.86 19.13 2.88 19.46 2.88 ;
        RECT  16.80 4.00 19.38 4.32 ;
        POLYGON  18.06 3.08 17.88 3.08 17.88 3.68 16.44 3.68 16.44 4.32
                 16.12 4.32 16.12 3.68 15.00 3.68 15.00 3.06 12.52 3.06
                 12.52 2.52 12.84 2.52 12.84 2.74 15.00 2.74 15.00 1.86
                 16.13 1.86 16.13 2.18 15.32 2.18 15.32 3.36 17.56 3.36
                 17.56 2.76 18.06 2.76 ;
        POLYGON  14.68 3.90 13.68 3.90 13.68 3.46 14.00 3.46 14.00 3.58
                 14.68 3.58 ;
        POLYGON  14.16 4.54 11.78 4.54 11.24 4.00 11.24 3.26 8.52 3.26
                 7.74 2.48 7.74 1.86 8.06 1.86 8.06 2.34 8.66 2.94 11.56 2.94
                 11.56 3.86 11.92 4.22 14.16 4.22 ;
        RECT  12.82 1.28 13.98 1.60 ;
        POLYGON  13.30 3.90 12.06 3.90 11.88 3.72 11.88 2.62 9.76 2.62
                 9.76 2.30 11.88 2.30 11.88 1.96 11.98 1.86 12.08 1.86
                 12.08 1.28 12.40 1.28 12.40 2.18 12.20 2.18 12.20 3.58
                 13.30 3.58 ;
        POLYGON  11.70 1.60 11.38 1.60 11.38 1.54 4.62 1.54 4.62 1.22
                 11.70 1.22 ;
        RECT  4.62 4.22 11.00 4.54 ;
        RECT  7.76 3.58 10.32 3.90 ;
        RECT  8.46 1.86 9.46 2.18 ;
        POLYGON  7.26 2.20 6.94 2.20 6.94 2.18 6.32 2.18 6.32 3.90 6.00 3.90
                 6.00 1.86 7.26 1.86 ;
        POLYGON  5.64 2.18 1.86 2.18 1.86 1.22 2.18 1.22 2.18 1.86 5.64 1.86 ;
        POLYGON  5.64 3.72 5.32 3.72 5.32 3.70 2.54 3.70 2.54 3.38 5.64 3.38 ;
        RECT  2.54 1.22 4.24 1.54 ;
        POLYGON  4.24 4.34 1.86 4.34 1.86 3.38 2.18 3.38 2.18 4.02 4.24 4.02 ;
        POLYGON  3.24 3.04 0.48 3.04 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.72 2.92 2.72
                 2.92 2.60 3.24 2.60 ;
    END
END sdffnrsq_2

MACRO sdffnrsq_1
    CLASS CORE ;
    FOREIGN sdffnrsq_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 28.80 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.96 3.04 15.84 3.04 15.84 2.72 16.64 2.72 16.64 2.50
                 16.96 2.50 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.62 4.56 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  28.00 2.40 27.74 2.40 27.74 3.28 27.59 3.28 27.59 4.54
                 27.27 4.54 27.27 2.96 27.42 2.96 27.42 1.54 27.27 1.54
                 27.27 1.22 27.74 1.22 27.74 2.08 28.00 2.08 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.52 3.04 6.80 3.04 6.80 2.60 7.20 2.60 7.20 2.72 7.52 2.72 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  23.16 2.62 23.52 3.26 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.95 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.76 1.12 2.40 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  28.80 0.90 26.09 0.90 26.09 1.52 25.77 1.52 25.77 0.90
                 23.01 0.90 23.01 1.53 22.69 1.53 22.69 0.90 1.33 0.90
                 1.33 1.12 1.01 1.12 1.01 0.90 0.00 0.90 0.00 -0.90 28.80 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  28.80 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.22 1.32 4.22
                 1.32 4.86 3.24 4.86 3.24 4.66 3.56 4.66 3.56 4.86 15.22 4.86
                 15.22 4.14 15.54 4.14 15.54 4.64 17.98 4.64 17.98 4.86
                 21.14 4.86 21.14 4.60 21.46 4.60 21.46 4.86 25.70 4.86
                 25.70 4.24 26.02 4.24 26.02 4.86 27.97 4.86 27.97 4.22
                 28.29 4.22 28.29 4.86 28.80 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  27.07 2.46 26.88 2.46 26.88 4.54 26.56 4.54 26.56 1.22
                 26.91 1.22 26.91 1.54 26.88 1.54 26.88 2.14 27.07 2.14 ;
        POLYGON  26.13 2.57 25.27 2.57 25.27 3.90 22.84 3.90 22.84 4.54
                 22.52 4.54 22.52 3.58 22.25 3.58 22.25 3.26 22.84 3.26
                 22.84 3.58 24.95 3.58 24.95 1.22 25.27 1.22 25.27 2.25
                 26.13 2.25 ;
        RECT  23.27 4.22 25.20 4.54 ;
        RECT  23.57 1.22 24.57 1.54 ;
        POLYGON  24.16 2.64 23.84 2.64 23.84 2.24 21.93 2.24 21.93 3.64
                 20.08 3.64 20.08 4.54 19.76 4.54 19.76 3.32 21.61 3.32
                 21.61 2.24 20.19 2.24 20.19 1.28 20.51 1.28 20.51 1.92
                 24.16 1.92 ;
        RECT  20.89 1.28 22.21 1.60 ;
        POLYGON  22.16 4.28 20.78 4.28 20.78 4.44 20.46 4.44 20.46 3.96
                 22.16 3.96 ;
        POLYGON  19.81 1.60 19.49 1.60 19.49 1.54 17.17 1.54 17.17 1.22
                 19.81 1.22 ;
        POLYGON  19.46 3.20 18.70 3.20 18.70 3.68 18.38 3.68 18.38 2.88
                 18.81 2.88 18.81 2.18 16.45 2.18 16.45 1.54 14.62 1.54
                 14.62 2.40 13.48 2.40 13.48 2.08 14.30 2.08 14.30 1.22
                 16.77 1.22 16.77 1.86 19.13 1.86 19.13 2.88 19.46 2.88 ;
        RECT  16.80 4.00 19.38 4.32 ;
        POLYGON  18.06 3.08 17.88 3.08 17.88 3.68 16.44 3.68 16.44 4.32
                 16.12 4.32 16.12 3.68 15.00 3.68 15.00 3.06 12.52 3.06
                 12.52 2.52 12.84 2.52 12.84 2.74 15.00 2.74 15.00 1.86
                 16.13 1.86 16.13 2.18 15.32 2.18 15.32 3.36 17.56 3.36
                 17.56 2.76 18.06 2.76 ;
        POLYGON  14.68 3.90 13.68 3.90 13.68 3.46 14.00 3.46 14.00 3.58
                 14.68 3.58 ;
        POLYGON  14.16 4.54 11.78 4.54 11.24 4.00 11.24 3.26 8.52 3.26
                 7.74 2.48 7.74 1.86 8.06 1.86 8.06 2.34 8.66 2.94 11.56 2.94
                 11.56 3.86 11.92 4.22 14.16 4.22 ;
        RECT  12.82 1.28 13.98 1.60 ;
        POLYGON  13.30 3.90 12.06 3.90 11.88 3.72 11.88 2.62 9.76 2.62
                 9.76 2.30 11.88 2.30 11.88 1.96 11.98 1.86 12.08 1.86
                 12.08 1.28 12.40 1.28 12.40 2.18 12.20 2.18 12.20 3.58
                 13.30 3.58 ;
        POLYGON  11.70 1.60 11.38 1.60 11.38 1.54 4.62 1.54 4.62 1.22
                 11.70 1.22 ;
        RECT  4.62 4.22 11.00 4.54 ;
        RECT  7.76 3.58 10.32 3.90 ;
        RECT  8.46 1.86 9.46 2.18 ;
        POLYGON  7.26 2.20 6.94 2.20 6.94 2.18 6.32 2.18 6.32 3.90 6.00 3.90
                 6.00 1.86 7.26 1.86 ;
        POLYGON  5.64 2.18 1.86 2.18 1.86 1.22 2.18 1.22 2.18 1.86 5.64 1.86 ;
        POLYGON  5.64 3.72 5.32 3.72 5.32 3.70 2.54 3.70 2.54 3.38 5.64 3.38 ;
        RECT  2.54 1.22 4.24 1.54 ;
        POLYGON  4.24 4.34 1.86 4.34 1.86 3.38 2.18 3.38 2.18 4.02 4.24 4.02 ;
        POLYGON  3.24 3.04 0.48 3.04 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.72 2.92 2.72
                 2.92 2.60 3.24 2.60 ;
    END
END sdffnrsq_1

MACRO sdffnrs_4
    CLASS CORE ;
    FOREIGN sdffnrs_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 32.00 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.96 3.04 15.84 3.04 15.84 2.72 16.64 2.72 16.64 2.50
                 16.96 2.50 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.62 4.56 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  29.52 3.25 27.75 3.25 27.75 2.93 28.96 2.93 28.96 2.72
                 29.20 2.72 29.20 1.87 27.27 1.87 27.27 1.55 29.52 1.55 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  31.84 4.53 29.84 4.53 29.84 4.21 31.52 4.21 31.52 1.90
                 29.84 1.90 29.84 1.58 31.84 1.58 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.52 3.04 6.80 3.04 6.80 2.60 7.20 2.60 7.20 2.72 7.52 2.72 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  23.16 2.62 23.52 3.26 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.95 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.76 1.12 2.40 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  32.00 0.90 30.86 0.90 30.86 1.23 30.54 1.23 30.54 0.90
                 28.29 0.90 28.29 1.23 27.97 1.23 27.97 0.90 25.97 0.90
                 25.97 1.52 25.65 1.52 25.65 0.90 23.01 0.90 23.01 1.53
                 22.69 1.53 22.69 0.90 1.32 0.90 1.32 1.12 1.00 1.12 1.00 0.90
                 0.00 0.90 0.00 -0.90 32.00 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  32.00 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.22 1.32 4.22
                 1.32 4.86 3.24 4.86 3.24 4.66 3.56 4.66 3.56 4.86 15.22 4.86
                 15.22 4.14 15.54 4.14 15.54 4.64 17.98 4.64 17.98 4.86
                 21.14 4.86 21.14 4.60 21.46 4.60 21.46 4.86 28.46 4.86
                 28.46 4.79 28.81 4.79 28.81 4.86 32.00 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  30.86 3.89 28.79 3.89 28.79 4.02 25.45 4.02 25.45 3.90
                 22.84 3.90 22.84 4.54 22.52 4.54 22.52 3.58 22.25 3.58
                 22.25 3.26 22.84 3.26 22.84 3.58 24.95 3.58 24.95 1.22
                 25.27 1.22 25.27 2.25 26.13 2.25 26.13 2.57 25.27 2.57
                 25.27 3.58 25.77 3.58 25.77 3.70 28.47 3.70 28.47 3.57
                 30.54 3.57 30.54 2.32 30.86 2.32 ;
        POLYGON  27.07 2.45 26.88 2.45 26.88 3.38 26.56 3.38 26.56 1.22
                 26.91 1.22 26.91 1.54 26.88 1.54 26.88 2.13 27.07 2.13 ;
        RECT  23.27 4.22 25.20 4.54 ;
        RECT  23.57 1.22 24.57 1.54 ;
        POLYGON  24.16 2.64 23.84 2.64 23.84 2.24 21.93 2.24 21.93 3.64
                 20.08 3.64 20.08 4.54 19.76 4.54 19.76 3.32 21.61 3.32
                 21.61 2.24 20.19 2.24 20.19 1.28 20.51 1.28 20.51 1.92
                 24.16 1.92 ;
        RECT  20.89 1.28 22.21 1.60 ;
        POLYGON  22.16 4.28 20.78 4.28 20.78 4.44 20.46 4.44 20.46 3.96
                 22.16 3.96 ;
        POLYGON  19.81 1.60 19.49 1.60 19.49 1.54 17.17 1.54 17.17 1.22
                 19.81 1.22 ;
        POLYGON  19.46 3.20 18.70 3.20 18.70 3.68 18.38 3.68 18.38 2.88
                 18.81 2.88 18.81 2.18 16.45 2.18 16.45 1.54 14.62 1.54
                 14.62 2.40 13.48 2.40 13.48 2.08 14.30 2.08 14.30 1.22
                 16.77 1.22 16.77 1.86 19.13 1.86 19.13 2.88 19.46 2.88 ;
        RECT  16.80 4.00 19.38 4.32 ;
        POLYGON  18.06 3.08 17.88 3.08 17.88 3.68 16.44 3.68 16.44 4.32
                 16.12 4.32 16.12 3.68 15.00 3.68 15.00 3.06 12.52 3.06
                 12.52 2.52 12.84 2.52 12.84 2.74 15.00 2.74 15.00 1.86
                 16.13 1.86 16.13 2.18 15.32 2.18 15.32 3.36 17.56 3.36
                 17.56 2.76 18.06 2.76 ;
        POLYGON  14.68 3.90 13.68 3.90 13.68 3.46 14.00 3.46 14.00 3.58
                 14.68 3.58 ;
        POLYGON  14.16 4.54 11.78 4.54 11.24 4.00 11.24 3.26 8.52 3.26
                 7.74 2.48 7.74 1.86 8.06 1.86 8.06 2.34 8.66 2.94 11.56 2.94
                 11.56 3.86 11.92 4.22 14.16 4.22 ;
        RECT  12.82 1.28 13.98 1.60 ;
        POLYGON  13.30 3.90 12.06 3.90 11.88 3.72 11.88 2.62 9.76 2.62
                 9.76 2.30 11.88 2.30 11.88 1.96 11.98 1.86 12.08 1.86
                 12.08 1.28 12.40 1.28 12.40 2.18 12.20 2.18 12.20 3.58
                 13.30 3.58 ;
        POLYGON  11.70 1.60 11.38 1.60 11.38 1.54 4.62 1.54 4.62 1.22
                 11.70 1.22 ;
        RECT  4.62 4.22 11.00 4.54 ;
        RECT  7.76 3.58 10.32 3.90 ;
        RECT  8.46 1.86 9.46 2.18 ;
        POLYGON  7.26 2.20 6.94 2.20 6.94 2.18 6.32 2.18 6.32 3.90 6.00 3.90
                 6.00 1.86 7.26 1.86 ;
        POLYGON  5.64 2.18 1.86 2.18 1.86 1.22 2.18 1.22 2.18 1.86 5.64 1.86 ;
        POLYGON  5.64 3.72 5.32 3.72 5.32 3.70 2.54 3.70 2.54 3.38 5.64 3.38 ;
        RECT  2.54 1.22 4.24 1.54 ;
        POLYGON  4.24 4.34 1.86 4.34 1.86 3.38 2.18 3.38 2.18 4.02 4.24 4.02 ;
        POLYGON  3.24 3.04 0.48 3.04 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.72 2.92 2.72
                 2.92 2.60 3.24 2.60 ;
    END
END sdffnrs_4

MACRO sdffnrs_2
    CLASS CORE ;
    FOREIGN sdffnrs_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 29.44 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.96 3.04 15.84 3.04 15.84 2.72 16.64 2.72 16.64 2.50
                 16.96 2.50 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.62 4.56 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.86  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  28.00 1.76 27.72 1.76 27.72 3.38 27.32 3.38 27.32 3.06
                 27.40 3.06 27.40 1.22 27.72 1.22 27.72 1.44 28.00 1.44 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  29.28 4.54 28.84 4.54 28.84 4.22 28.96 4.22 28.96 1.54
                 28.84 1.54 28.84 1.22 29.28 1.22 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.52 3.04 6.80 3.04 6.80 2.60 7.20 2.60 7.20 2.72 7.52 2.72 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  23.16 2.62 23.52 3.26 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.95 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.76 1.12 2.40 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  29.44 0.90 25.97 0.90 25.97 1.52 25.65 1.52 25.65 0.90
                 23.01 0.90 23.01 1.53 22.69 1.53 22.69 0.90 1.32 0.90
                 1.32 1.12 1.00 1.12 1.00 0.90 0.00 0.90 0.00 -0.90 29.44 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  29.44 6.66 0.00 6.66 0.00 4.86 1.03 4.86 1.03 4.22 1.35 4.22
                 1.35 4.86 3.24 4.86 3.24 4.66 3.56 4.66 3.56 4.86 15.22 4.86
                 15.22 4.14 15.54 4.14 15.54 4.64 17.98 4.64 17.98 4.86
                 21.14 4.86 21.14 4.60 21.46 4.60 21.46 4.86 29.44 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  28.58 4.02 25.45 4.02 25.45 3.90 22.84 3.90 22.84 4.54
                 22.52 4.54 22.52 3.58 22.25 3.58 22.25 3.26 22.84 3.26
                 22.84 3.58 24.95 3.58 24.95 1.22 25.27 1.22 25.27 2.25
                 26.13 2.25 26.13 2.57 25.27 2.57 25.27 3.58 25.77 3.58
                 25.77 3.70 28.26 3.70 28.26 2.12 28.58 2.12 ;
        POLYGON  27.07 2.46 26.88 2.46 26.88 3.06 26.92 3.06 26.92 3.38
                 26.56 3.38 26.56 1.22 26.91 1.22 26.91 1.54 26.88 1.54
                 26.88 2.14 27.07 2.14 ;
        RECT  23.27 4.22 25.20 4.54 ;
        RECT  23.57 1.22 24.57 1.54 ;
        POLYGON  24.16 2.64 23.84 2.64 23.84 2.24 21.93 2.24 21.93 3.64
                 20.08 3.64 20.08 4.54 19.76 4.54 19.76 3.32 21.61 3.32
                 21.61 2.24 20.19 2.24 20.19 1.28 20.51 1.28 20.51 1.92
                 24.16 1.92 ;
        RECT  20.89 1.28 22.21 1.60 ;
        POLYGON  22.16 4.28 20.78 4.28 20.78 4.44 20.46 4.44 20.46 3.96
                 22.16 3.96 ;
        POLYGON  19.81 1.60 19.49 1.60 19.49 1.54 17.17 1.54 17.17 1.22
                 19.81 1.22 ;
        POLYGON  19.46 3.20 18.70 3.20 18.70 3.68 18.38 3.68 18.38 2.88
                 18.81 2.88 18.81 2.18 16.45 2.18 16.45 1.54 14.62 1.54
                 14.62 2.40 13.48 2.40 13.48 2.08 14.30 2.08 14.30 1.22
                 16.77 1.22 16.77 1.86 19.13 1.86 19.13 2.88 19.46 2.88 ;
        RECT  16.80 4.00 19.38 4.32 ;
        POLYGON  18.06 3.08 17.88 3.08 17.88 3.68 16.44 3.68 16.44 4.32
                 16.12 4.32 16.12 3.68 15.00 3.68 15.00 3.06 12.52 3.06
                 12.52 2.52 12.84 2.52 12.84 2.74 15.00 2.74 15.00 1.86
                 16.13 1.86 16.13 2.18 15.32 2.18 15.32 3.36 17.56 3.36
                 17.56 2.76 18.06 2.76 ;
        POLYGON  14.68 3.90 13.68 3.90 13.68 3.46 14.00 3.46 14.00 3.58
                 14.68 3.58 ;
        POLYGON  14.16 4.54 11.78 4.54 11.24 4.00 11.24 3.26 8.52 3.26
                 7.74 2.48 7.74 1.86 8.06 1.86 8.06 2.34 8.66 2.94 11.56 2.94
                 11.56 3.86 11.92 4.22 14.16 4.22 ;
        RECT  12.82 1.28 13.98 1.60 ;
        POLYGON  13.30 3.90 12.06 3.90 11.88 3.72 11.88 2.62 9.76 2.62
                 9.76 2.30 11.88 2.30 11.88 1.96 11.98 1.86 12.08 1.86
                 12.08 1.28 12.40 1.28 12.40 2.18 12.20 2.18 12.20 3.58
                 13.30 3.58 ;
        POLYGON  11.70 1.60 11.38 1.60 11.38 1.54 4.62 1.54 4.62 1.22
                 11.70 1.22 ;
        RECT  4.62 4.22 11.00 4.54 ;
        RECT  7.76 3.58 10.32 3.90 ;
        RECT  8.46 1.86 9.46 2.18 ;
        POLYGON  7.26 2.20 6.94 2.20 6.94 2.18 6.32 2.18 6.32 3.90 6.00 3.90
                 6.00 1.86 7.26 1.86 ;
        POLYGON  5.64 2.18 1.86 2.18 1.86 1.22 2.18 1.22 2.18 1.86 5.64 1.86 ;
        POLYGON  5.64 3.72 5.32 3.72 5.32 3.70 2.54 3.70 2.54 3.38 5.64 3.38 ;
        RECT  2.54 1.22 4.24 1.54 ;
        POLYGON  4.24 4.34 1.86 4.34 1.86 3.38 2.18 3.38 2.18 4.02 4.24 4.02 ;
        POLYGON  3.24 3.04 0.48 3.04 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.72 2.92 2.72
                 2.92 2.60 3.24 2.60 ;
    END
END sdffnrs_2

MACRO sdffnrs_1
    CLASS CORE ;
    FOREIGN sdffnrs_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 29.44 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.96 3.04 15.84 3.04 15.84 2.72 16.64 2.72 16.64 2.50
                 16.96 2.50 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.62 4.56 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.43  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  28.00 1.76 27.72 1.76 27.72 3.38 27.32 3.38 27.32 3.06
                 27.40 3.06 27.40 1.22 27.72 1.22 27.72 1.44 28.00 1.44 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  29.28 4.54 28.84 4.54 28.84 4.22 28.96 4.22 28.96 1.54
                 28.84 1.54 28.84 1.22 29.28 1.22 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.52 3.04 6.80 3.04 6.80 2.60 7.20 2.60 7.20 2.72 7.52 2.72 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  23.16 2.62 23.52 3.26 ;
        END
    END sb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.67  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.95 2.62 5.60 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.76 1.12 2.40 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  29.44 0.90 26.10 0.90 26.10 1.52 25.78 1.52 25.78 0.90
                 23.01 0.90 23.01 1.53 22.69 1.53 22.69 0.90 1.32 0.90
                 1.32 1.12 1.00 1.12 1.00 0.90 0.00 0.90 0.00 -0.90 29.44 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  29.44 6.66 0.00 6.66 0.00 4.86 0.99 4.86 0.99 4.22 1.31 4.22
                 1.31 4.86 3.24 4.86 3.24 4.66 3.56 4.66 3.56 4.86 15.22 4.86
                 15.22 4.14 15.54 4.14 15.54 4.64 17.98 4.64 17.98 4.86
                 21.14 4.86 21.14 4.60 21.46 4.60 21.46 4.86 28.12 4.86
                 28.12 4.58 28.44 4.58 28.44 4.86 29.44 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  28.58 4.02 25.45 4.02 25.45 3.90 22.84 3.90 22.84 4.54
                 22.52 4.54 22.52 3.58 22.25 3.58 22.25 3.26 22.84 3.26
                 22.84 3.58 24.95 3.58 24.95 1.22 25.27 1.22 25.27 2.25
                 26.13 2.25 26.13 2.57 25.27 2.57 25.27 3.58 25.77 3.58
                 25.77 3.70 28.26 3.70 28.26 2.12 28.58 2.12 ;
        POLYGON  27.07 2.46 26.88 2.46 26.88 3.06 26.92 3.06 26.92 3.38
                 26.56 3.38 26.56 1.22 26.91 1.22 26.91 1.54 26.88 1.54
                 26.88 2.14 27.07 2.14 ;
        RECT  23.27 4.22 25.20 4.54 ;
        RECT  23.57 1.22 24.57 1.54 ;
        POLYGON  24.16 2.64 23.84 2.64 23.84 2.24 21.93 2.24 21.93 3.64
                 20.08 3.64 20.08 4.54 19.76 4.54 19.76 3.32 21.61 3.32
                 21.61 2.24 20.19 2.24 20.19 1.28 20.51 1.28 20.51 1.92
                 24.16 1.92 ;
        RECT  20.89 1.28 22.21 1.60 ;
        POLYGON  22.16 4.28 20.78 4.28 20.78 4.44 20.46 4.44 20.46 3.96
                 22.16 3.96 ;
        POLYGON  19.81 1.60 19.49 1.60 19.49 1.54 17.17 1.54 17.17 1.22
                 19.81 1.22 ;
        POLYGON  19.46 3.20 18.70 3.20 18.70 3.68 18.38 3.68 18.38 2.88
                 18.81 2.88 18.81 2.18 16.45 2.18 16.45 1.54 14.62 1.54
                 14.62 2.40 13.48 2.40 13.48 2.08 14.30 2.08 14.30 1.22
                 16.77 1.22 16.77 1.86 19.13 1.86 19.13 2.88 19.46 2.88 ;
        RECT  16.80 4.00 19.38 4.32 ;
        POLYGON  18.06 3.08 17.88 3.08 17.88 3.68 16.44 3.68 16.44 4.32
                 16.12 4.32 16.12 3.68 15.00 3.68 15.00 3.06 12.52 3.06
                 12.52 2.52 12.84 2.52 12.84 2.74 15.00 2.74 15.00 1.86
                 16.13 1.86 16.13 2.18 15.32 2.18 15.32 3.36 17.56 3.36
                 17.56 2.76 18.06 2.76 ;
        POLYGON  14.68 3.90 13.68 3.90 13.68 3.46 14.00 3.46 14.00 3.58
                 14.68 3.58 ;
        POLYGON  14.16 4.54 11.78 4.54 11.24 4.00 11.24 3.26 8.52 3.26
                 7.74 2.48 7.74 1.86 8.06 1.86 8.06 2.34 8.66 2.94 11.56 2.94
                 11.56 3.86 11.92 4.22 14.16 4.22 ;
        RECT  12.82 1.28 13.98 1.60 ;
        POLYGON  13.30 3.90 12.06 3.90 11.88 3.72 11.88 2.62 9.76 2.62
                 9.76 2.30 11.88 2.30 11.88 1.96 11.98 1.86 12.08 1.86
                 12.08 1.28 12.40 1.28 12.40 2.18 12.20 2.18 12.20 3.58
                 13.30 3.58 ;
        POLYGON  11.70 1.60 11.38 1.60 11.38 1.54 4.62 1.54 4.62 1.22
                 11.70 1.22 ;
        RECT  4.62 4.22 11.00 4.54 ;
        RECT  7.76 3.58 10.32 3.90 ;
        RECT  8.46 1.86 9.46 2.18 ;
        POLYGON  7.26 2.20 6.94 2.20 6.94 2.18 6.32 2.18 6.32 3.90 6.00 3.90
                 6.00 1.86 7.26 1.86 ;
        POLYGON  5.64 2.18 1.86 2.18 1.86 1.22 2.18 1.22 2.18 1.86 5.64 1.86 ;
        POLYGON  5.64 3.72 5.32 3.72 5.32 3.70 2.54 3.70 2.54 3.38 5.64 3.38 ;
        RECT  2.54 1.22 4.24 1.54 ;
        POLYGON  4.24 4.34 1.86 4.34 1.86 3.38 2.18 3.38 2.18 4.02 4.24 4.02 ;
        POLYGON  3.24 3.04 0.48 3.04 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.72 2.92 2.72
                 2.92 2.60 3.24 2.60 ;
    END
END sdffnrs_1

MACRO sdffnrqb_4
    CLASS CORE ;
    FOREIGN sdffnrqb_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 26.88 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  13.52 2.72 14.18 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.65 5.28 3.04 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  26.72 3.04 26.48 3.04 26.48 4.54 24.76 4.54 24.76 4.22
                 26.16 4.22 26.16 1.54 24.76 1.54 24.76 1.22 26.48 1.22
                 26.48 2.72 26.72 2.72 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.44  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  8.48 2.08 8.94 2.62 ;
        END
    END rb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.60 2.65 6.34 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.65 3.04 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  26.88 0.90 23.46 0.90 23.46 1.54 23.14 1.54 23.14 0.90
                 14.04 0.90 14.04 1.54 13.72 1.54 13.72 0.90 1.88 0.90
                 1.88 1.71 0.88 1.71 0.88 0.90 0.00 0.90 0.00 -0.90 26.88 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  26.88 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 21.76 4.86 21.76 4.12 22.08 4.12 22.08 4.86
                 23.26 4.86 23.26 4.22 23.58 4.22 23.58 4.86 26.88 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  25.75 2.46 24.40 2.46 24.40 4.54 24.08 4.54 24.08 3.16
                 21.80 3.16 21.80 2.84 24.08 2.84 24.08 1.54 23.84 1.54
                 23.84 1.22 24.40 1.22 24.40 2.14 25.75 2.14 ;
        POLYGON  23.64 2.52 21.48 2.52 21.48 3.48 22.76 3.48 22.76 4.54
                 22.44 4.54 22.44 3.80 20.14 3.80 19.90 4.04 19.90 4.54
                 19.58 4.54 19.58 3.90 20.00 3.48 21.16 3.48 21.16 2.52
                 20.44 2.52 19.68 1.76 19.68 1.22 20.00 1.22 20.00 1.62
                 20.58 2.20 23.64 2.20 ;
        RECT  21.76 1.22 22.76 1.54 ;
        RECT  20.38 1.22 21.38 1.54 ;
        RECT  20.28 4.12 21.38 4.44 ;
        POLYGON  19.42 3.24 18.76 3.90 17.66 3.90 17.66 4.54 13.86 4.54
                 13.86 4.05 13.71 3.90 12.54 3.90 12.54 3.26 11.16 3.26
                 11.16 2.94 12.86 2.94 12.86 3.58 13.85 3.58 14.18 3.91
                 14.18 4.22 17.34 4.22 17.34 3.58 18.62 3.58 19.10 3.10
                 19.10 2.50 18.78 2.18 16.06 2.18 16.06 1.86 18.92 1.86
                 19.42 2.36 ;
        RECT  18.30 1.22 19.30 1.54 ;
        RECT  18.20 4.22 19.20 4.54 ;
        POLYGON  18.78 2.96 17.02 2.96 17.02 3.90 14.50 3.90 14.50 2.18
                 11.48 2.18 11.48 2.56 11.16 2.56 11.16 1.86 14.82 1.86
                 14.82 3.58 16.70 3.58 16.70 2.64 18.78 2.64 ;
        POLYGON  17.92 1.54 15.74 1.54 15.74 2.54 16.28 2.54 16.28 2.86
                 15.42 2.86 15.42 1.22 17.92 1.22 ;
        POLYGON  13.54 4.54 9.88 4.54 9.88 3.90 6.86 3.90 6.86 2.68 7.22 2.32
                 7.22 1.87 7.54 1.87 7.54 2.46 7.18 2.82 7.18 3.58 10.20 3.58
                 10.20 4.22 13.54 4.22 ;
        RECT  12.34 1.22 13.34 1.54 ;
        RECT  11.22 3.58 12.22 3.90 ;
        RECT  10.96 1.22 11.96 1.54 ;
        POLYGON  10.84 3.90 10.52 3.90 10.52 3.26 7.52 3.26 7.52 2.94
                 10.26 2.94 10.26 1.22 10.58 1.22 10.58 2.94 10.84 2.94 ;
        RECT  5.84 1.22 9.88 1.54 ;
        RECT  5.48 4.22 9.56 4.54 ;
        RECT  2.94 1.87 6.86 2.19 ;
        RECT  4.10 3.58 6.50 3.90 ;
        RECT  4.34 1.23 5.34 1.55 ;
        RECT  2.70 4.22 5.10 4.54 ;
        POLYGON  4.26 2.97 3.78 2.97 3.78 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 1.87 0.50 1.87 0.50 3.58 3.46 3.58 3.46 2.65 4.26 2.65 ;
        POLYGON  3.96 1.55 2.58 1.55 2.58 2.19 2.26 2.19 2.26 1.23 3.96 1.23 ;
    END
END sdffnrqb_4

MACRO sdffnrqb_2
    CLASS CORE ;
    FOREIGN sdffnrqb_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 26.24 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  13.52 2.72 14.18 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.65 5.28 3.04 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.69  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  26.08 1.76 25.90 1.76 25.90 4.54 25.47 4.54 25.47 4.22
                 25.58 4.22 25.58 1.54 25.46 1.54 25.46 1.22 25.90 1.22
                 25.90 1.44 26.08 1.44 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.44  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  8.48 2.08 8.94 2.62 ;
        END
    END rb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.60 2.65 6.34 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.65 3.04 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  26.24 0.90 23.46 0.90 23.46 1.54 23.14 1.54 23.14 0.90
                 14.04 0.90 14.04 1.54 13.72 1.54 13.72 0.90 1.88 0.90
                 1.88 1.71 0.88 1.71 0.88 0.90 0.00 0.90 0.00 -0.90 26.24 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  26.24 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 21.76 4.86 21.76 4.12 22.08 4.12 22.08 4.86
                 23.26 4.86 23.26 4.22 23.58 4.22 23.58 4.86 26.24 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  25.26 2.44 25.02 2.44 25.02 3.07 25.01 3.07 25.01 3.16
                 24.28 3.16 24.28 4.22 24.44 4.22 24.44 4.54 23.96 4.54
                 23.96 3.16 21.80 3.16 21.80 2.84 23.96 2.84 23.96 1.54
                 23.84 1.54 23.84 1.22 24.28 1.22 24.28 2.84 24.70 2.84
                 24.70 2.12 25.26 2.12 ;
        POLYGON  23.64 2.52 21.48 2.52 21.48 3.48 22.76 3.48 22.76 4.54
                 22.44 4.54 22.44 3.80 20.14 3.80 19.90 4.04 19.90 4.54
                 19.58 4.54 19.58 3.90 20.00 3.48 21.16 3.48 21.16 2.52
                 20.44 2.52 19.68 1.76 19.68 1.22 20.00 1.22 20.00 1.62
                 20.58 2.20 23.64 2.20 ;
        RECT  21.76 1.22 22.76 1.54 ;
        RECT  20.38 1.22 21.38 1.54 ;
        RECT  20.28 4.12 21.38 4.44 ;
        POLYGON  19.42 3.24 18.76 3.90 17.66 3.90 17.66 4.54 13.86 4.54
                 13.86 4.05 13.71 3.90 12.54 3.90 12.54 3.26 11.16 3.26
                 11.16 2.94 12.86 2.94 12.86 3.58 13.85 3.58 14.18 3.91
                 14.18 4.22 17.34 4.22 17.34 3.58 18.62 3.58 19.10 3.10
                 19.10 2.50 18.78 2.18 16.06 2.18 16.06 1.86 18.92 1.86
                 19.42 2.36 ;
        RECT  18.30 1.22 19.30 1.54 ;
        RECT  18.20 4.22 19.20 4.54 ;
        POLYGON  18.78 2.96 17.02 2.96 17.02 3.90 14.50 3.90 14.50 2.18
                 11.48 2.18 11.48 2.56 11.16 2.56 11.16 1.86 14.82 1.86
                 14.82 3.58 16.70 3.58 16.70 2.64 18.78 2.64 ;
        POLYGON  17.92 1.54 15.74 1.54 15.74 2.54 16.28 2.54 16.28 2.86
                 15.42 2.86 15.42 1.22 17.92 1.22 ;
        POLYGON  13.54 4.54 9.88 4.54 9.88 3.90 6.86 3.90 6.86 2.68 7.22 2.32
                 7.22 1.87 7.54 1.87 7.54 2.46 7.18 2.82 7.18 3.58 10.20 3.58
                 10.20 4.22 13.54 4.22 ;
        RECT  12.34 1.22 13.34 1.54 ;
        RECT  11.22 3.58 12.22 3.90 ;
        RECT  10.96 1.22 11.96 1.54 ;
        POLYGON  10.84 3.90 10.52 3.90 10.52 3.26 7.52 3.26 7.52 2.94
                 10.26 2.94 10.26 1.22 10.58 1.22 10.58 2.94 10.84 2.94 ;
        RECT  5.84 1.22 9.88 1.54 ;
        RECT  5.48 4.22 9.56 4.54 ;
        RECT  2.94 1.87 6.86 2.19 ;
        RECT  4.10 3.58 6.50 3.90 ;
        RECT  4.34 1.23 5.34 1.55 ;
        RECT  2.70 4.22 5.10 4.54 ;
        POLYGON  4.26 2.97 3.78 2.97 3.78 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 1.87 0.50 1.87 0.50 3.58 3.46 3.58 3.46 2.65 4.26 2.65 ;
        POLYGON  3.96 1.55 2.58 1.55 2.58 2.19 2.26 2.19 2.26 1.23 3.96 1.23 ;
    END
END sdffnrqb_2

MACRO sdffnrqb_1
    CLASS CORE ;
    FOREIGN sdffnrqb_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 26.24 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  13.52 2.72 14.18 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.65 5.28 3.04 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.23  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  26.08 1.76 25.90 1.76 25.90 4.54 25.47 4.54 25.47 4.22
                 25.58 4.22 25.58 1.54 25.46 1.54 25.46 1.22 25.90 1.22
                 25.90 1.44 26.08 1.44 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.44  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  8.48 2.08 8.94 2.62 ;
        END
    END rb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.60 2.65 6.34 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.65 3.04 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  26.24 0.90 23.46 0.90 23.46 1.54 23.14 1.54 23.14 0.90
                 14.04 0.90 14.04 1.54 13.72 1.54 13.72 0.90 1.88 0.90
                 1.88 1.71 0.88 1.71 0.88 0.90 0.00 0.90 0.00 -0.90 26.24 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  26.24 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 21.76 4.86 21.76 4.12 22.08 4.12 22.08 4.86
                 23.26 4.86 23.26 4.22 23.58 4.22 23.58 4.86 26.24 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  25.26 3.39 25.02 3.39 25.02 3.96 23.96 3.96 23.96 3.16
                 21.80 3.16 21.80 2.84 23.96 2.84 23.96 1.54 23.84 1.54
                 23.84 1.22 24.28 1.22 24.28 3.64 24.70 3.64 24.70 3.07
                 25.26 3.07 ;
        POLYGON  23.64 2.52 21.48 2.52 21.48 3.48 22.76 3.48 22.76 4.54
                 22.44 4.54 22.44 3.80 20.14 3.80 19.90 4.04 19.90 4.54
                 19.58 4.54 19.58 3.90 20.00 3.48 21.16 3.48 21.16 2.52
                 20.44 2.52 19.68 1.76 19.68 1.22 20.00 1.22 20.00 1.62
                 20.58 2.20 23.64 2.20 ;
        RECT  21.76 1.22 22.76 1.54 ;
        RECT  20.38 1.22 21.38 1.54 ;
        RECT  20.28 4.12 21.38 4.44 ;
        POLYGON  19.42 3.24 18.76 3.90 17.66 3.90 17.66 4.54 13.86 4.54
                 13.86 4.05 13.71 3.90 12.54 3.90 12.54 3.26 11.16 3.26
                 11.16 2.94 12.86 2.94 12.86 3.58 13.85 3.58 14.18 3.91
                 14.18 4.22 17.34 4.22 17.34 3.58 18.62 3.58 19.10 3.10
                 19.10 2.50 18.78 2.18 16.06 2.18 16.06 1.86 18.92 1.86
                 19.42 2.36 ;
        RECT  18.30 1.22 19.30 1.54 ;
        RECT  18.20 4.22 19.20 4.54 ;
        POLYGON  18.78 2.96 17.02 2.96 17.02 3.90 14.50 3.90 14.50 2.18
                 11.48 2.18 11.48 2.56 11.16 2.56 11.16 1.86 14.82 1.86
                 14.82 3.58 16.70 3.58 16.70 2.64 18.78 2.64 ;
        POLYGON  17.92 1.54 15.74 1.54 15.74 2.54 16.28 2.54 16.28 2.86
                 15.42 2.86 15.42 1.22 17.92 1.22 ;
        POLYGON  13.54 4.54 9.88 4.54 9.88 3.90 6.86 3.90 6.86 2.68 7.22 2.32
                 7.22 1.87 7.54 1.87 7.54 2.46 7.18 2.82 7.18 3.58 10.20 3.58
                 10.20 4.22 13.54 4.22 ;
        RECT  12.34 1.22 13.34 1.54 ;
        RECT  11.22 3.58 12.22 3.90 ;
        RECT  10.96 1.22 11.96 1.54 ;
        POLYGON  10.84 3.90 10.52 3.90 10.52 3.26 7.52 3.26 7.52 2.94
                 10.26 2.94 10.26 1.22 10.58 1.22 10.58 2.94 10.84 2.94 ;
        RECT  5.84 1.22 9.88 1.54 ;
        RECT  5.48 4.22 9.56 4.54 ;
        RECT  2.94 1.87 6.86 2.19 ;
        RECT  4.10 3.58 6.50 3.90 ;
        RECT  4.34 1.23 5.34 1.55 ;
        RECT  2.70 4.22 5.10 4.54 ;
        POLYGON  4.26 2.97 3.78 2.97 3.78 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 1.87 0.50 1.87 0.50 3.58 3.46 3.58 3.46 2.65 4.26 2.65 ;
        POLYGON  3.96 1.55 2.58 1.55 2.58 2.19 2.26 2.19 2.26 1.23 3.96 1.23 ;
    END
END sdffnrqb_1

MACRO sdffnrq_4
    CLASS CORE ;
    FOREIGN sdffnrq_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 26.88 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  13.52 2.72 14.18 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.65 5.28 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  26.48 4.54 26.16 4.54 26.16 3.04 25.08 3.04 25.08 4.54
                 24.76 4.54 24.76 1.22 25.08 1.22 25.08 2.72 26.16 2.72
                 26.16 1.22 26.48 1.22 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.44  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  8.48 2.08 8.94 2.62 ;
        END
    END rb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.60 2.65 6.34 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.65 3.04 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  26.88 0.90 25.78 0.90 25.78 1.54 25.46 1.54 25.46 0.90
                 23.46 0.90 23.46 1.54 23.14 1.54 23.14 0.90 14.04 0.90
                 14.04 1.54 13.72 1.54 13.72 0.90 1.88 0.90 1.88 1.71 0.88 1.71
                 0.88 0.90 0.00 0.90 0.00 -0.90 26.88 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  26.88 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 21.76 4.86 21.76 4.22 22.08 4.22 22.08 4.86
                 23.26 4.86 23.26 4.22 23.58 4.22 23.58 4.86 25.46 4.86
                 25.46 3.58 25.78 3.58 25.78 4.86 26.88 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  24.40 4.54 24.08 4.54 24.08 3.16 21.80 3.16 21.80 2.84
                 24.08 2.84 24.08 1.54 23.84 1.54 23.84 1.22 24.40 1.22 ;
        POLYGON  23.64 2.52 21.48 2.52 21.48 3.48 22.76 3.48 22.76 4.54
                 22.44 4.54 22.44 3.80 20.14 3.80 19.90 4.04 19.90 4.54
                 19.58 4.54 19.58 3.90 20.00 3.48 21.16 3.48 21.16 2.52
                 20.44 2.52 19.68 1.76 19.68 1.22 20.00 1.22 20.00 1.62
                 20.58 2.20 23.64 2.20 ;
        RECT  21.76 1.22 22.76 1.54 ;
        RECT  20.38 1.22 21.38 1.54 ;
        RECT  20.28 4.22 21.38 4.54 ;
        POLYGON  19.42 3.24 18.76 3.90 17.66 3.90 17.66 4.54 13.86 4.54
                 13.86 4.05 13.71 3.90 12.54 3.90 12.54 3.26 11.16 3.26
                 11.16 2.94 12.86 2.94 12.86 3.58 13.85 3.58 14.18 3.91
                 14.18 4.22 17.34 4.22 17.34 3.58 18.62 3.58 19.10 3.10
                 19.10 2.50 18.78 2.18 16.06 2.18 16.06 1.86 18.92 1.86
                 19.42 2.36 ;
        RECT  18.30 1.22 19.30 1.54 ;
        RECT  18.20 4.22 19.20 4.54 ;
        POLYGON  18.78 2.96 17.02 2.96 17.02 3.90 14.50 3.90 14.50 2.18
                 11.48 2.18 11.48 2.56 11.16 2.56 11.16 1.86 14.82 1.86
                 14.82 3.58 16.70 3.58 16.70 2.64 18.78 2.64 ;
        POLYGON  17.92 1.54 15.74 1.54 15.74 2.54 16.28 2.54 16.28 2.86
                 15.42 2.86 15.42 1.22 17.92 1.22 ;
        POLYGON  13.54 4.54 9.88 4.54 9.88 3.90 6.86 3.90 6.86 2.68 7.22 2.32
                 7.22 1.87 7.54 1.87 7.54 2.46 7.18 2.82 7.18 3.58 10.20 3.58
                 10.20 4.22 13.54 4.22 ;
        RECT  12.34 1.22 13.34 1.54 ;
        RECT  11.22 3.58 12.22 3.90 ;
        RECT  10.96 1.22 11.96 1.54 ;
        POLYGON  10.84 3.90 10.52 3.90 10.52 3.26 7.52 3.26 7.52 2.94
                 10.26 2.94 10.26 1.22 10.58 1.22 10.58 2.94 10.84 2.94 ;
        RECT  5.84 1.22 9.88 1.54 ;
        RECT  5.48 4.22 9.56 4.54 ;
        RECT  2.94 1.87 6.86 2.19 ;
        RECT  4.10 3.58 6.50 3.90 ;
        RECT  4.34 1.23 5.34 1.55 ;
        RECT  2.70 4.22 5.10 4.54 ;
        POLYGON  4.26 2.97 3.78 2.97 3.78 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 1.87 0.50 1.87 0.50 3.58 3.46 3.58 3.46 2.65 4.26 2.65 ;
        POLYGON  3.96 1.55 2.58 1.55 2.58 2.19 2.26 2.19 2.26 1.23 3.96 1.23 ;
    END
END sdffnrq_4

MACRO sdffnrq_2
    CLASS CORE ;
    FOREIGN sdffnrq_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 26.24 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  13.52 2.72 14.18 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.65 5.28 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  25.44 3.04 25.08 3.04 25.08 4.54 24.76 4.54 24.76 1.22
                 25.08 1.22 25.08 2.72 25.44 2.72 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.44  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  8.48 2.08 8.94 2.62 ;
        END
    END rb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.60 2.65 6.34 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.65 3.04 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  26.24 0.90 25.78 0.90 25.78 1.54 25.46 1.54 25.46 0.90
                 23.46 0.90 23.46 1.54 23.14 1.54 23.14 0.90 14.04 0.90
                 14.04 1.54 13.72 1.54 13.72 0.90 1.88 0.90 1.88 1.71 0.88 1.71
                 0.88 0.90 0.00 0.90 0.00 -0.90 26.24 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  26.24 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 21.76 4.86 21.76 4.12 22.08 4.12 22.08 4.86
                 23.26 4.86 23.26 4.22 23.58 4.22 23.58 4.86 25.46 4.86
                 25.46 3.58 25.78 3.58 25.78 4.86 26.24 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  24.40 4.54 24.08 4.54 24.08 3.16 21.80 3.16 21.80 2.84
                 24.08 2.84 24.08 1.54 23.84 1.54 23.84 1.22 24.40 1.22 ;
        POLYGON  23.64 2.52 21.48 2.52 21.48 3.48 22.76 3.48 22.76 4.54
                 22.44 4.54 22.44 3.80 20.14 3.80 19.90 4.04 19.90 4.54
                 19.58 4.54 19.58 3.90 20.00 3.48 21.16 3.48 21.16 2.52
                 20.44 2.52 19.68 1.76 19.68 1.22 20.00 1.22 20.00 1.62
                 20.58 2.20 23.64 2.20 ;
        RECT  21.76 1.22 22.76 1.54 ;
        RECT  20.38 1.22 21.38 1.54 ;
        RECT  20.28 4.12 21.38 4.44 ;
        POLYGON  19.42 3.24 18.76 3.90 17.66 3.90 17.66 4.54 13.86 4.54
                 13.86 4.05 13.71 3.90 12.54 3.90 12.54 3.26 11.16 3.26
                 11.16 2.94 12.86 2.94 12.86 3.58 13.85 3.58 14.18 3.91
                 14.18 4.22 17.34 4.22 17.34 3.58 18.62 3.58 19.10 3.10
                 19.10 2.50 18.78 2.18 16.06 2.18 16.06 1.86 18.92 1.86
                 19.42 2.36 ;
        RECT  18.30 1.22 19.30 1.54 ;
        RECT  18.20 4.22 19.20 4.54 ;
        POLYGON  18.78 2.96 17.02 2.96 17.02 3.90 14.50 3.90 14.50 2.18
                 11.48 2.18 11.48 2.56 11.16 2.56 11.16 1.86 14.82 1.86
                 14.82 3.58 16.70 3.58 16.70 2.64 18.78 2.64 ;
        POLYGON  17.92 1.54 15.74 1.54 15.74 2.54 16.28 2.54 16.28 2.86
                 15.42 2.86 15.42 1.22 17.92 1.22 ;
        POLYGON  13.54 4.54 9.88 4.54 9.88 3.90 6.86 3.90 6.86 2.68 7.22 2.32
                 7.22 1.87 7.54 1.87 7.54 2.46 7.18 2.82 7.18 3.58 10.20 3.58
                 10.20 4.22 13.54 4.22 ;
        RECT  12.34 1.22 13.34 1.54 ;
        RECT  11.22 3.58 12.22 3.90 ;
        RECT  10.96 1.22 11.96 1.54 ;
        POLYGON  10.84 3.90 10.52 3.90 10.52 3.26 7.52 3.26 7.52 2.94
                 10.26 2.94 10.26 1.22 10.58 1.22 10.58 2.94 10.84 2.94 ;
        RECT  5.84 1.22 9.88 1.54 ;
        RECT  5.48 4.22 9.56 4.54 ;
        RECT  2.94 1.87 6.86 2.19 ;
        RECT  4.10 3.58 6.50 3.90 ;
        RECT  4.34 1.23 5.34 1.55 ;
        RECT  2.70 4.22 5.10 4.54 ;
        POLYGON  4.26 2.97 3.78 2.97 3.78 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 1.87 0.50 1.87 0.50 3.58 3.46 3.58 3.46 2.65 4.26 2.65 ;
        POLYGON  3.96 1.55 2.58 1.55 2.58 2.19 2.26 2.19 2.26 1.23 3.96 1.23 ;
    END
END sdffnrq_2

MACRO sdffnrq_1
    CLASS CORE ;
    FOREIGN sdffnrq_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 26.24 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  13.52 2.72 14.18 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.65 5.28 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  25.44 3.04 25.08 3.04 25.08 4.44 24.76 4.44 24.76 1.22
                 25.08 1.22 25.08 2.72 25.44 2.72 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.44  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  8.48 2.08 8.94 2.62 ;
        END
    END rb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.60 2.65 6.34 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.65 3.04 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  26.24 0.90 25.78 0.90 25.78 1.24 25.46 1.24 25.46 0.90
                 23.46 0.90 23.46 1.54 23.14 1.54 23.14 0.90 14.04 0.90
                 14.04 1.54 13.72 1.54 13.72 0.90 1.88 0.90 1.88 1.71 0.88 1.71
                 0.88 0.90 0.00 0.90 0.00 -0.90 26.24 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  26.24 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 21.76 4.86 21.76 4.12 22.08 4.12 22.08 4.86
                 23.26 4.86 23.26 4.12 23.58 4.12 23.58 4.86 25.46 4.86
                 25.46 4.12 25.78 4.12 25.78 4.86 26.24 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  24.40 4.44 24.08 4.44 24.08 3.16 21.80 3.16 21.80 2.84
                 24.08 2.84 24.08 1.54 23.84 1.54 23.84 1.22 24.40 1.22 ;
        POLYGON  23.64 2.52 21.48 2.52 21.48 3.48 22.76 3.48 22.76 4.44
                 22.44 4.44 22.44 3.80 20.14 3.80 19.90 4.04 19.90 4.54
                 19.58 4.54 19.58 3.90 20.00 3.48 21.16 3.48 21.16 2.52
                 20.44 2.52 19.68 1.76 19.68 1.22 20.00 1.22 20.00 1.62
                 20.58 2.20 23.64 2.20 ;
        RECT  21.76 1.22 22.76 1.54 ;
        RECT  20.38 1.22 21.38 1.54 ;
        RECT  20.28 4.12 21.38 4.44 ;
        POLYGON  19.42 3.24 18.76 3.90 17.66 3.90 17.66 4.54 13.86 4.54
                 13.86 4.05 13.71 3.90 12.54 3.90 12.54 3.26 11.16 3.26
                 11.16 2.94 12.86 2.94 12.86 3.58 13.85 3.58 14.18 3.91
                 14.18 4.22 17.34 4.22 17.34 3.58 18.62 3.58 19.10 3.10
                 19.10 2.50 18.78 2.18 16.06 2.18 16.06 1.86 18.92 1.86
                 19.42 2.36 ;
        RECT  18.30 1.22 19.30 1.54 ;
        RECT  18.20 4.22 19.20 4.54 ;
        POLYGON  18.78 2.96 17.02 2.96 17.02 3.90 14.50 3.90 14.50 2.18
                 11.48 2.18 11.48 2.56 11.16 2.56 11.16 1.86 14.82 1.86
                 14.82 3.58 16.70 3.58 16.70 2.64 18.78 2.64 ;
        POLYGON  17.92 1.54 15.74 1.54 15.74 2.54 16.28 2.54 16.28 2.86
                 15.42 2.86 15.42 1.22 17.92 1.22 ;
        POLYGON  13.54 4.54 9.88 4.54 9.88 3.90 6.86 3.90 6.86 2.68 7.22 2.32
                 7.22 1.87 7.54 1.87 7.54 2.46 7.18 2.82 7.18 3.58 10.20 3.58
                 10.20 4.22 13.54 4.22 ;
        RECT  12.34 1.22 13.34 1.54 ;
        RECT  11.22 3.58 12.22 3.90 ;
        RECT  10.96 1.22 11.96 1.54 ;
        POLYGON  10.84 3.90 10.52 3.90 10.52 3.26 7.52 3.26 7.52 2.94
                 10.26 2.94 10.26 1.22 10.58 1.22 10.58 2.94 10.84 2.94 ;
        RECT  5.84 1.22 9.88 1.54 ;
        RECT  5.48 4.22 9.56 4.54 ;
        RECT  2.94 1.87 6.86 2.19 ;
        RECT  4.10 3.58 6.50 3.90 ;
        RECT  4.34 1.23 5.34 1.55 ;
        RECT  2.70 4.22 5.10 4.54 ;
        POLYGON  4.26 2.97 3.78 2.97 3.78 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 1.87 0.50 1.87 0.50 3.58 3.46 3.58 3.46 2.65 4.26 2.65 ;
        POLYGON  3.96 1.55 2.58 1.55 2.58 2.19 2.26 2.19 2.26 1.23 3.96 1.23 ;
    END
END sdffnrq_1

MACRO sdffnr_4
    CLASS CORE ;
    FOREIGN sdffnr_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 28.80 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  13.52 2.72 14.18 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.65 5.28 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.35  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  26.49 3.26 24.72 3.26 24.72 1.22 26.48 1.22 26.48 1.54
                 25.04 1.54 25.04 2.72 25.44 2.72 25.44 2.94 26.49 2.94 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  28.64 3.04 28.57 3.04 28.57 4.54 26.85 4.54 26.85 4.22
                 28.25 4.22 28.25 1.54 26.85 1.54 26.85 1.22 28.57 1.22
                 28.57 2.72 28.64 2.72 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.44  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  8.48 2.08 8.94 2.62 ;
        END
    END rb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.60 2.65 6.34 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.65 3.04 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  28.80 0.90 23.46 0.90 23.46 1.54 23.14 1.54 23.14 0.90
                 14.04 0.90 14.04 1.54 13.72 1.54 13.72 0.90 1.88 0.90
                 1.88 1.71 0.88 1.71 0.88 0.90 0.00 0.90 0.00 -0.90 28.80 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  28.80 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 21.76 4.86 21.76 4.12 22.08 4.12 22.08 4.86
                 23.26 4.86 23.26 4.22 23.58 4.22 23.58 4.86 25.46 4.86
                 25.46 4.22 25.78 4.22 25.78 4.86 28.80 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  27.88 2.46 27.13 2.46 27.13 3.90 24.40 3.90 24.40 4.54
                 24.08 4.54 24.08 3.16 21.80 3.16 21.80 2.84 24.08 2.84
                 24.08 1.54 23.84 1.54 23.84 1.22 24.40 1.22 24.40 3.58
                 26.81 3.58 26.81 2.14 27.88 2.14 ;
        POLYGON  23.64 2.52 21.48 2.52 21.48 3.48 22.76 3.48 22.76 4.54
                 22.44 4.54 22.44 3.80 20.14 3.80 19.90 4.04 19.90 4.54
                 19.58 4.54 19.58 3.90 20.00 3.48 21.16 3.48 21.16 2.52
                 20.44 2.52 19.68 1.76 19.68 1.22 20.00 1.22 20.00 1.62
                 20.58 2.20 23.64 2.20 ;
        RECT  21.76 1.22 22.76 1.54 ;
        RECT  20.38 1.22 21.38 1.54 ;
        RECT  20.28 4.12 21.38 4.44 ;
        POLYGON  19.42 3.24 18.76 3.90 17.66 3.90 17.66 4.54 13.86 4.54
                 13.86 4.05 13.71 3.90 12.54 3.90 12.54 3.26 11.16 3.26
                 11.16 2.94 12.86 2.94 12.86 3.58 13.85 3.58 14.18 3.91
                 14.18 4.22 17.34 4.22 17.34 3.58 18.62 3.58 19.10 3.10
                 19.10 2.50 18.78 2.18 16.06 2.18 16.06 1.86 18.92 1.86
                 19.42 2.36 ;
        RECT  18.30 1.22 19.30 1.54 ;
        RECT  18.20 4.22 19.20 4.54 ;
        POLYGON  18.78 2.96 17.02 2.96 17.02 3.90 14.50 3.90 14.50 2.18
                 11.48 2.18 11.48 2.56 11.16 2.56 11.16 1.86 14.82 1.86
                 14.82 3.58 16.70 3.58 16.70 2.64 18.78 2.64 ;
        POLYGON  17.92 1.54 15.74 1.54 15.74 2.54 16.28 2.54 16.28 2.86
                 15.42 2.86 15.42 1.22 17.92 1.22 ;
        POLYGON  13.54 4.54 9.88 4.54 9.88 3.90 6.86 3.90 6.86 2.68 7.22 2.32
                 7.22 1.87 7.54 1.87 7.54 2.46 7.18 2.82 7.18 3.58 10.20 3.58
                 10.20 4.22 13.54 4.22 ;
        RECT  12.34 1.22 13.34 1.54 ;
        RECT  11.22 3.58 12.22 3.90 ;
        RECT  10.96 1.22 11.96 1.54 ;
        POLYGON  10.84 3.90 10.52 3.90 10.52 3.26 7.52 3.26 7.52 2.94
                 10.26 2.94 10.26 1.22 10.58 1.22 10.58 2.94 10.84 2.94 ;
        RECT  5.84 1.22 9.88 1.54 ;
        RECT  5.48 4.22 9.56 4.54 ;
        RECT  2.94 1.87 6.86 2.19 ;
        RECT  4.10 3.58 6.50 3.90 ;
        RECT  4.34 1.23 5.34 1.55 ;
        RECT  2.70 4.22 5.10 4.54 ;
        POLYGON  4.26 2.97 3.78 2.97 3.78 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 1.87 0.50 1.87 0.50 3.58 3.46 3.58 3.46 2.65 4.26 2.65 ;
        POLYGON  3.96 1.55 2.58 1.55 2.58 2.19 2.26 2.19 2.26 1.23 3.96 1.23 ;
    END
END sdffnr_4

MACRO sdffnr_2
    CLASS CORE ;
    FOREIGN sdffnr_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 26.88 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  13.52 2.72 14.18 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.65 5.28 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  25.44 1.76 25.04 1.76 25.04 3.58 25.08 3.58 25.08 3.90
                 24.72 3.90 24.72 1.22 25.44 1.22 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.69  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  26.72 1.76 26.60 1.76 26.60 4.54 26.17 4.54 26.17 4.22
                 26.28 4.22 26.28 1.54 26.16 1.54 26.16 1.22 26.60 1.22
                 26.60 1.44 26.72 1.44 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.44  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  8.48 2.08 8.94 2.62 ;
        END
    END rb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.60 2.65 6.34 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.65 3.04 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  26.88 0.90 23.46 0.90 23.46 1.54 23.14 1.54 23.14 0.90
                 14.04 0.90 14.04 1.54 13.72 1.54 13.72 0.90 1.88 0.90
                 1.88 1.71 0.88 1.71 0.88 0.90 0.00 0.90 0.00 -0.90 26.88 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  26.88 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 21.76 4.86 21.76 4.12 22.08 4.12 22.08 4.86
                 23.26 4.86 23.26 4.22 23.58 4.22 23.58 4.86 26.88 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  25.96 2.44 25.72 2.44 25.72 4.54 23.96 4.54 23.96 3.16
                 21.80 3.16 21.80 2.84 23.96 2.84 23.96 1.54 23.84 1.54
                 23.84 1.22 24.28 1.22 24.28 4.22 25.40 4.22 25.40 2.12
                 25.96 2.12 ;
        POLYGON  23.64 2.52 21.48 2.52 21.48 3.48 22.76 3.48 22.76 4.54
                 22.44 4.54 22.44 3.80 20.14 3.80 19.90 4.04 19.90 4.54
                 19.58 4.54 19.58 3.90 20.00 3.48 21.16 3.48 21.16 2.52
                 20.44 2.52 19.68 1.76 19.68 1.22 20.00 1.22 20.00 1.62
                 20.58 2.20 23.64 2.20 ;
        RECT  21.76 1.22 22.76 1.54 ;
        RECT  20.38 1.22 21.38 1.54 ;
        RECT  20.28 4.12 21.38 4.44 ;
        POLYGON  19.42 3.24 18.76 3.90 17.66 3.90 17.66 4.54 13.86 4.54
                 13.86 4.05 13.71 3.90 12.54 3.90 12.54 3.26 11.16 3.26
                 11.16 2.94 12.86 2.94 12.86 3.58 13.85 3.58 14.18 3.91
                 14.18 4.22 17.34 4.22 17.34 3.58 18.62 3.58 19.10 3.10
                 19.10 2.50 18.78 2.18 16.06 2.18 16.06 1.86 18.92 1.86
                 19.42 2.36 ;
        RECT  18.30 1.22 19.30 1.54 ;
        RECT  18.20 4.22 19.20 4.54 ;
        POLYGON  18.78 2.96 17.02 2.96 17.02 3.90 14.50 3.90 14.50 2.18
                 11.48 2.18 11.48 2.56 11.16 2.56 11.16 1.86 14.82 1.86
                 14.82 3.58 16.70 3.58 16.70 2.64 18.78 2.64 ;
        POLYGON  17.92 1.54 15.74 1.54 15.74 2.54 16.28 2.54 16.28 2.86
                 15.42 2.86 15.42 1.22 17.92 1.22 ;
        POLYGON  13.54 4.54 9.88 4.54 9.88 3.90 6.86 3.90 6.86 2.68 7.22 2.32
                 7.22 1.87 7.54 1.87 7.54 2.46 7.18 2.82 7.18 3.58 10.20 3.58
                 10.20 4.22 13.54 4.22 ;
        RECT  12.34 1.22 13.34 1.54 ;
        RECT  11.22 3.58 12.22 3.90 ;
        RECT  10.96 1.22 11.96 1.54 ;
        POLYGON  10.84 3.90 10.52 3.90 10.52 3.26 7.52 3.26 7.52 2.94
                 10.26 2.94 10.26 1.22 10.58 1.22 10.58 2.94 10.84 2.94 ;
        RECT  5.84 1.22 9.88 1.54 ;
        RECT  5.48 4.22 9.56 4.54 ;
        RECT  2.94 1.87 6.86 2.19 ;
        RECT  4.10 3.58 6.50 3.90 ;
        RECT  4.34 1.23 5.34 1.55 ;
        RECT  2.70 4.22 5.10 4.54 ;
        POLYGON  4.26 2.97 3.78 2.97 3.78 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 1.87 0.50 1.87 0.50 3.58 3.46 3.58 3.46 2.65 4.26 2.65 ;
        POLYGON  3.96 1.55 2.58 1.55 2.58 2.19 2.26 2.19 2.26 1.23 3.96 1.23 ;
    END
END sdffnr_2

MACRO sdffnr_1
    CLASS CORE ;
    FOREIGN sdffnr_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 26.88 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  13.52 2.72 14.18 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.65 5.28 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.21  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  25.44 1.76 25.04 1.76 25.04 3.58 25.08 3.58 25.08 3.90
                 24.72 3.90 24.72 1.22 25.44 1.22 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.23  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  26.72 1.76 26.60 1.76 26.60 4.54 26.17 4.54 26.17 4.22
                 26.28 4.22 26.28 1.54 26.16 1.54 26.16 1.22 26.60 1.22
                 26.60 1.44 26.72 1.44 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.44  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  8.48 2.08 8.94 2.62 ;
        END
    END rb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.60 2.65 6.34 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.65 3.04 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  26.88 0.90 23.46 0.90 23.46 1.54 23.14 1.54 23.14 0.90
                 14.04 0.90 14.04 1.54 13.72 1.54 13.72 0.90 1.88 0.90
                 1.88 1.71 0.88 1.71 0.88 0.90 0.00 0.90 0.00 -0.90 26.88 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  26.88 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 21.76 4.86 21.76 4.12 22.08 4.12 22.08 4.86
                 23.26 4.86 23.26 4.22 23.58 4.22 23.58 4.86 26.88 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  25.96 2.44 25.72 2.44 25.72 4.54 23.96 4.54 23.96 3.16
                 21.80 3.16 21.80 2.84 23.96 2.84 23.96 1.54 23.84 1.54
                 23.84 1.22 24.28 1.22 24.28 4.22 25.40 4.22 25.40 2.12
                 25.96 2.12 ;
        POLYGON  23.64 2.52 21.48 2.52 21.48 3.48 22.76 3.48 22.76 4.54
                 22.44 4.54 22.44 3.80 20.14 3.80 19.90 4.04 19.90 4.54
                 19.58 4.54 19.58 3.90 20.00 3.48 21.16 3.48 21.16 2.52
                 20.44 2.52 19.68 1.76 19.68 1.22 20.00 1.22 20.00 1.62
                 20.58 2.20 23.64 2.20 ;
        RECT  21.76 1.22 22.76 1.54 ;
        RECT  20.38 1.22 21.38 1.54 ;
        RECT  20.28 4.12 21.38 4.44 ;
        POLYGON  19.42 3.24 18.76 3.90 17.66 3.90 17.66 4.54 13.86 4.54
                 13.86 4.05 13.71 3.90 12.54 3.90 12.54 3.26 11.16 3.26
                 11.16 2.94 12.86 2.94 12.86 3.58 13.85 3.58 14.18 3.91
                 14.18 4.22 17.34 4.22 17.34 3.58 18.62 3.58 19.10 3.10
                 19.10 2.50 18.78 2.18 16.06 2.18 16.06 1.86 18.92 1.86
                 19.42 2.36 ;
        RECT  18.30 1.22 19.30 1.54 ;
        RECT  18.20 4.22 19.20 4.54 ;
        POLYGON  18.78 2.96 17.02 2.96 17.02 3.90 14.50 3.90 14.50 2.18
                 11.48 2.18 11.48 2.56 11.16 2.56 11.16 1.86 14.82 1.86
                 14.82 3.58 16.70 3.58 16.70 2.64 18.78 2.64 ;
        POLYGON  17.92 1.54 15.74 1.54 15.74 2.54 16.28 2.54 16.28 2.86
                 15.42 2.86 15.42 1.22 17.92 1.22 ;
        POLYGON  13.54 4.54 9.88 4.54 9.88 3.90 6.86 3.90 6.86 2.68 7.22 2.32
                 7.22 1.87 7.54 1.87 7.54 2.46 7.18 2.82 7.18 3.58 10.20 3.58
                 10.20 4.22 13.54 4.22 ;
        RECT  12.34 1.22 13.34 1.54 ;
        RECT  11.22 3.58 12.22 3.90 ;
        RECT  10.96 1.22 11.96 1.54 ;
        POLYGON  10.84 3.90 10.52 3.90 10.52 3.26 7.52 3.26 7.52 2.94
                 10.26 2.94 10.26 1.22 10.58 1.22 10.58 2.94 10.84 2.94 ;
        RECT  5.84 1.22 9.88 1.54 ;
        RECT  5.48 4.22 9.56 4.54 ;
        RECT  2.94 1.87 6.86 2.19 ;
        RECT  4.10 3.58 6.50 3.90 ;
        RECT  4.34 1.23 5.34 1.55 ;
        RECT  2.70 4.22 5.10 4.54 ;
        POLYGON  4.26 2.97 3.78 2.97 3.78 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 1.87 0.50 1.87 0.50 3.58 3.46 3.58 3.46 2.65 4.26 2.65 ;
        POLYGON  3.96 1.55 2.58 1.55 2.58 2.19 2.26 2.19 2.26 1.23 3.96 1.23 ;
    END
END sdffnr_1

MACRO sdffnqb_4
    CLASS CORE ;
    FOREIGN sdffnqb_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  13.63 3.46 12.64 3.46 12.64 3.68 12.32 3.68 12.32 3.14
                 13.63 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.68 2.66 4.32 3.04 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.96 4.53 19.09 4.53 19.09 4.21 20.64 4.21 20.64 1.90
                 19.09 1.90 19.09 1.58 20.96 1.58 ;
        END
    END qb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.66 5.28 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.66 1.76 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 0.90 20.11 0.90 20.11 1.23 19.55 1.23 19.55 0.90
                 17.79 0.90 17.79 1.14 17.47 1.14 17.47 0.90 10.30 0.90
                 10.30 1.48 9.98 1.48 9.98 0.90 2.58 0.90 2.58 1.54 2.26 1.54
                 2.26 0.90 1.20 0.90 1.20 1.86 0.88 1.86 0.88 0.90 0.00 0.90
                 0.00 -0.90 21.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 10.54 4.86 10.54 3.74 10.86 3.74 10.86 4.86
                 17.53 4.86 17.53 3.96 17.85 3.96 17.85 4.86 21.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.11 2.66 18.49 2.66 18.49 3.53 18.76 3.53 18.76 3.85
                 18.17 3.85 18.17 3.18 17.19 3.18 17.19 2.86 18.17 2.86
                 18.17 1.22 18.49 1.22 18.49 2.34 20.11 2.34 ;
        POLYGON  17.85 2.47 17.53 2.47 17.53 2.28 15.63 2.28 15.63 4.54
                 15.31 4.54 15.31 2.28 14.87 1.84 14.87 1.22 15.19 1.22
                 15.19 1.70 15.45 1.96 17.85 1.96 ;
        RECT  16.09 3.96 17.09 4.28 ;
        RECT  15.69 1.22 16.99 1.54 ;
        RECT  11.97 4.22 14.93 4.54 ;
        POLYGON  14.77 3.90 13.93 3.90 13.93 3.58 14.45 3.58 14.45 2.34
                 14.29 2.18 11.26 2.18 11.26 1.86 14.43 1.86 14.77 2.20 ;
        RECT  11.73 1.22 14.37 1.54 ;
        POLYGON  14.13 2.86 13.81 2.86 13.81 2.82 11.69 2.82 11.69 3.90
                 11.37 3.90 11.37 2.82 9.27 2.82 9.27 3.13 8.95 3.13 8.95 2.50
                 10.62 2.50 10.62 1.22 11.00 1.22 11.00 1.54 10.94 1.54
                 10.94 2.50 14.13 2.50 ;
        RECT  9.01 3.46 10.05 3.78 ;
        POLYGON  9.69 4.54 8.30 4.54 7.66 3.90 5.72 3.90 5.72 1.86 6.04 1.86
                 6.04 3.58 7.80 3.58 8.44 4.22 9.69 4.22 ;
        RECT  8.60 1.22 9.60 1.54 ;
        POLYGON  8.63 3.63 8.31 3.63 8.31 3.26 6.38 3.26 6.38 2.94 7.90 2.94
                 7.90 1.22 8.22 1.22 8.22 2.94 8.63 2.94 ;
        RECT  4.34 1.22 7.52 1.54 ;
        RECT  4.34 4.22 7.52 4.54 ;
        POLYGON  5.36 2.18 1.56 2.18 1.56 1.22 1.88 1.22 1.88 1.86 5.36 1.86 ;
        RECT  2.96 3.58 5.36 3.90 ;
        RECT  2.96 1.22 3.96 1.54 ;
        RECT  1.56 4.22 3.96 4.54 ;
        POLYGON  2.74 2.98 2.40 2.98 2.40 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 1.86 0.50 1.86 0.50 3.58 2.08 3.58 2.08 2.66 2.74 2.66 ;
    END
END sdffnqb_4

MACRO sdffnqb_2
    CLASS CORE ;
    FOREIGN sdffnqb_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 20.48 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  13.63 3.46 12.64 3.46 12.64 3.68 12.32 3.68 12.32 3.14
                 13.63 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.68 2.66 4.32 3.04 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.32 3.04 20.11 3.04 20.11 4.54 19.79 4.54 19.79 3.04
                 19.55 3.04 19.55 1.64 19.87 1.64 19.87 2.72 20.32 2.72 ;
        END
    END qb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.66 5.28 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.66 1.76 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 0.90 19.17 0.90 19.17 1.96 18.85 1.96 18.85 0.90
                 17.79 0.90 17.79 1.14 17.47 1.14 17.47 0.90 10.30 0.90
                 10.30 1.48 9.98 1.48 9.98 0.90 2.58 0.90 2.58 1.54 2.26 1.54
                 2.26 0.90 1.20 0.90 1.20 1.86 0.88 1.86 0.88 0.90 0.00 0.90
                 0.00 -0.90 20.48 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 10.54 4.86 10.54 3.74 10.86 3.74 10.86 4.86
                 17.53 4.86 17.53 3.96 17.85 3.96 17.85 4.86 19.09 4.86
                 19.09 4.22 19.41 4.22 19.41 4.86 20.48 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  19.23 2.94 18.49 2.94 18.49 4.22 18.73 4.22 18.73 4.54
                 18.17 4.54 18.17 3.18 17.19 3.18 17.19 2.86 18.17 2.86
                 18.17 1.22 18.49 1.22 18.49 2.62 19.23 2.62 ;
        POLYGON  17.85 2.47 17.53 2.47 17.53 2.28 15.63 2.28 15.63 4.54
                 15.31 4.54 15.31 2.28 14.87 1.84 14.87 1.22 15.19 1.22
                 15.19 1.70 15.45 1.96 17.85 1.96 ;
        RECT  16.09 3.96 17.09 4.28 ;
        RECT  15.69 1.22 16.99 1.54 ;
        RECT  11.97 4.22 14.93 4.54 ;
        POLYGON  14.77 3.90 13.93 3.90 13.93 3.58 14.45 3.58 14.45 2.34
                 14.29 2.18 11.26 2.18 11.26 1.86 14.43 1.86 14.77 2.20 ;
        RECT  11.73 1.22 14.37 1.54 ;
        POLYGON  14.13 2.86 13.81 2.86 13.81 2.82 11.69 2.82 11.69 3.90
                 11.37 3.90 11.37 2.82 9.27 2.82 9.27 3.13 8.95 3.13 8.95 2.50
                 10.62 2.50 10.62 1.22 11.00 1.22 11.00 1.54 10.94 1.54
                 10.94 2.50 14.13 2.50 ;
        RECT  9.01 3.46 10.05 3.78 ;
        POLYGON  9.69 4.54 8.30 4.54 7.66 3.90 5.72 3.90 5.72 1.86 6.04 1.86
                 6.04 3.58 7.80 3.58 8.44 4.22 9.69 4.22 ;
        RECT  8.60 1.22 9.60 1.54 ;
        POLYGON  8.63 3.63 8.31 3.63 8.31 3.26 6.38 3.26 6.38 2.94 7.90 2.94
                 7.90 1.22 8.22 1.22 8.22 2.94 8.63 2.94 ;
        RECT  4.34 1.22 7.52 1.54 ;
        RECT  4.34 4.22 7.52 4.54 ;
        POLYGON  5.36 2.18 1.56 2.18 1.56 1.22 1.88 1.22 1.88 1.86 5.36 1.86 ;
        RECT  2.96 3.58 5.36 3.90 ;
        RECT  2.96 1.22 3.96 1.54 ;
        RECT  1.56 4.22 3.96 4.54 ;
        POLYGON  2.74 2.98 2.40 2.98 2.40 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 1.86 0.50 1.86 0.50 3.58 2.08 3.58 2.08 2.66 2.74 2.66 ;
    END
END sdffnqb_2

MACRO sdffnqb_1
    CLASS CORE ;
    FOREIGN sdffnqb_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 20.48 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  13.63 3.46 12.64 3.46 12.64 3.68 12.32 3.68 12.32 3.14
                 13.63 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.68 2.66 4.32 3.04 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.32 4.54 19.88 4.54 19.88 4.22 20.00 4.22 20.00 1.54
                 19.55 1.54 19.55 1.22 20.32 1.22 ;
        END
    END qb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.66 5.28 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.66 1.76 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 0.90 19.17 0.90 19.17 1.54 18.85 1.54 18.85 0.90
                 17.79 0.90 17.79 1.54 17.47 1.54 17.47 0.90 10.30 0.90
                 10.30 1.48 9.98 1.48 9.98 0.90 2.58 0.90 2.58 1.54 2.26 1.54
                 2.26 0.90 1.20 0.90 1.20 1.86 0.88 1.86 0.88 0.90 0.00 0.90
                 0.00 -0.90 20.48 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 10.54 4.86 10.54 3.74 10.86 3.74 10.86 4.86
                 17.53 4.86 17.53 3.96 17.85 3.96 17.85 4.86 20.48 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  19.62 2.46 18.49 2.46 18.49 4.22 18.78 4.22 18.78 4.54
                 18.17 4.54 18.17 3.18 17.19 3.18 17.19 2.86 18.17 2.86
                 18.17 1.22 18.49 1.22 18.49 2.14 19.62 2.14 ;
        POLYGON  17.85 2.47 17.53 2.47 17.53 2.28 15.63 2.28 15.63 4.54
                 15.31 4.54 15.31 2.28 14.87 1.84 14.87 1.22 15.19 1.22
                 15.19 1.70 15.45 1.96 17.85 1.96 ;
        RECT  16.09 3.96 17.09 4.28 ;
        RECT  15.69 1.22 16.99 1.54 ;
        RECT  11.97 4.22 14.93 4.54 ;
        POLYGON  14.77 3.90 13.93 3.90 13.93 3.58 14.45 3.58 14.45 2.34
                 14.29 2.18 11.26 2.18 11.26 1.86 14.43 1.86 14.77 2.20 ;
        RECT  11.73 1.22 14.37 1.54 ;
        POLYGON  14.13 2.86 13.81 2.86 13.81 2.82 11.69 2.82 11.69 3.90
                 11.37 3.90 11.37 2.82 9.27 2.82 9.27 3.13 8.95 3.13 8.95 2.50
                 10.62 2.50 10.62 1.22 11.00 1.22 11.00 1.54 10.94 1.54
                 10.94 2.50 14.13 2.50 ;
        RECT  9.01 3.46 10.05 3.78 ;
        POLYGON  9.69 4.54 8.30 4.54 7.66 3.90 5.72 3.90 5.72 1.86 6.04 1.86
                 6.04 3.58 7.80 3.58 8.44 4.22 9.69 4.22 ;
        RECT  8.60 1.22 9.60 1.54 ;
        POLYGON  8.63 3.63 8.31 3.63 8.31 3.26 6.38 3.26 6.38 2.94 7.90 2.94
                 7.90 1.22 8.22 1.22 8.22 2.94 8.63 2.94 ;
        RECT  4.34 1.22 7.52 1.54 ;
        RECT  4.34 4.22 7.52 4.54 ;
        POLYGON  5.36 2.18 1.56 2.18 1.56 1.22 1.88 1.22 1.88 1.86 5.36 1.86 ;
        RECT  2.96 3.58 5.36 3.90 ;
        RECT  2.96 1.22 3.96 1.54 ;
        RECT  1.56 4.22 3.96 4.54 ;
        POLYGON  2.74 2.98 2.40 2.98 2.40 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 1.86 0.50 1.86 0.50 3.58 2.08 3.58 2.08 2.66 2.74 2.66 ;
    END
END sdffnqb_1

MACRO sdffnq_4
    CLASS CORE ;
    FOREIGN sdffnq_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  13.63 3.46 12.64 3.46 12.64 3.68 12.32 3.68 12.32 3.14
                 13.63 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.68 2.66 4.32 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.81 4.54 20.49 4.54 20.49 3.04 19.41 3.04 19.41 4.54
                 19.09 4.54 19.09 3.04 18.85 3.04 18.85 1.22 19.17 1.22
                 19.17 2.72 20.25 2.72 20.25 1.22 20.57 1.22 20.57 2.72
                 20.81 2.72 ;
        END
    END q
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.66 5.28 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.66 1.76 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 0.90 19.87 0.90 19.87 1.54 19.55 1.54 19.55 0.90
                 17.79 0.90 17.79 1.14 17.47 1.14 17.47 0.90 10.30 0.90
                 10.30 1.48 9.98 1.48 9.98 0.90 2.58 0.90 2.58 1.54 2.26 1.54
                 2.26 0.90 1.20 0.90 1.20 1.86 0.88 1.86 0.88 0.90 0.00 0.90
                 0.00 -0.90 21.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 10.54 4.86 10.54 3.74 10.86 3.74 10.86 4.86
                 17.53 4.86 17.53 3.96 17.85 3.96 17.85 4.86 19.79 4.86
                 19.79 3.58 20.11 3.58 20.11 4.86 21.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  18.73 4.54 18.17 4.54 18.17 3.18 17.19 3.18 17.19 2.86
                 18.17 2.86 18.17 1.22 18.49 1.22 18.49 4.22 18.73 4.22 ;
        POLYGON  17.85 2.47 17.53 2.47 17.53 2.28 15.63 2.28 15.63 4.54
                 15.31 4.54 15.31 2.28 14.87 1.84 14.87 1.22 15.19 1.22
                 15.19 1.70 15.45 1.96 17.85 1.96 ;
        RECT  16.09 3.96 17.09 4.28 ;
        RECT  15.69 1.22 16.99 1.54 ;
        RECT  11.97 4.22 14.93 4.54 ;
        POLYGON  14.77 3.90 13.93 3.90 13.93 3.58 14.45 3.58 14.45 2.34
                 14.29 2.18 11.26 2.18 11.26 1.86 14.43 1.86 14.77 2.20 ;
        RECT  11.73 1.22 14.37 1.54 ;
        POLYGON  14.13 2.86 13.81 2.86 13.81 2.82 11.69 2.82 11.69 3.90
                 11.37 3.90 11.37 2.82 9.27 2.82 9.27 3.13 8.95 3.13 8.95 2.50
                 10.62 2.50 10.62 1.22 11.00 1.22 11.00 1.54 10.94 1.54
                 10.94 2.50 14.13 2.50 ;
        RECT  9.01 3.46 10.05 3.78 ;
        POLYGON  9.69 4.54 8.30 4.54 7.66 3.90 5.72 3.90 5.72 1.86 6.04 1.86
                 6.04 3.58 7.80 3.58 8.44 4.22 9.69 4.22 ;
        RECT  8.60 1.22 9.60 1.54 ;
        POLYGON  8.63 3.63 8.31 3.63 8.31 3.26 6.38 3.26 6.38 2.94 7.90 2.94
                 7.90 1.22 8.22 1.22 8.22 2.94 8.63 2.94 ;
        RECT  4.34 1.22 7.52 1.54 ;
        RECT  4.34 4.22 7.52 4.54 ;
        POLYGON  5.36 2.18 1.56 2.18 1.56 1.22 1.88 1.22 1.88 1.86 5.36 1.86 ;
        RECT  2.96 3.58 5.36 3.90 ;
        RECT  2.96 1.22 3.96 1.54 ;
        RECT  1.56 4.22 3.96 4.54 ;
        POLYGON  2.74 2.98 2.40 2.98 2.40 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 1.86 0.50 1.86 0.50 3.58 2.08 3.58 2.08 2.66 2.74 2.66 ;
    END
END sdffnq_4

MACRO sdffnq_2
    CLASS CORE ;
    FOREIGN sdffnq_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 20.48 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  13.63 3.46 12.64 3.46 12.64 3.68 12.32 3.68 12.32 3.14
                 13.63 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.68 2.66 4.32 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.32 3.04 20.11 3.04 20.11 4.54 19.79 4.54 19.79 3.04
                 19.55 3.04 19.55 1.64 19.87 1.64 19.87 2.72 20.32 2.72 ;
        END
    END q
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.66 5.28 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.66 1.76 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 0.90 19.17 0.90 19.17 1.96 18.85 1.96 18.85 0.90
                 17.79 0.90 17.79 1.14 17.47 1.14 17.47 0.90 10.30 0.90
                 10.30 1.48 9.98 1.48 9.98 0.90 2.58 0.90 2.58 1.54 2.26 1.54
                 2.26 0.90 1.20 0.90 1.20 1.86 0.88 1.86 0.88 0.90 0.00 0.90
                 0.00 -0.90 20.48 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 10.54 4.86 10.54 3.74 10.86 3.74 10.86 4.86
                 17.53 4.86 17.53 3.96 17.85 3.96 17.85 4.86 19.09 4.86
                 19.09 4.22 19.41 4.22 19.41 4.86 20.48 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  18.73 4.54 18.17 4.54 18.17 3.18 17.19 3.18 17.19 2.86
                 18.17 2.86 18.17 1.22 18.49 1.22 18.49 4.22 18.73 4.22 ;
        POLYGON  17.85 2.47 17.53 2.47 17.53 2.28 15.63 2.28 15.63 4.54
                 15.31 4.54 15.31 2.28 14.87 1.84 14.87 1.22 15.19 1.22
                 15.19 1.70 15.45 1.96 17.85 1.96 ;
        RECT  16.09 3.96 17.09 4.28 ;
        RECT  15.69 1.22 16.99 1.54 ;
        RECT  11.97 4.22 14.93 4.54 ;
        POLYGON  14.77 3.90 13.93 3.90 13.93 3.58 14.45 3.58 14.45 2.34
                 14.29 2.18 11.26 2.18 11.26 1.86 14.43 1.86 14.77 2.20 ;
        RECT  11.73 1.22 14.37 1.54 ;
        POLYGON  14.13 2.86 13.81 2.86 13.81 2.82 11.69 2.82 11.69 3.90
                 11.37 3.90 11.37 2.82 9.27 2.82 9.27 3.13 8.95 3.13 8.95 2.50
                 10.62 2.50 10.62 1.22 11.00 1.22 11.00 1.54 10.94 1.54
                 10.94 2.50 14.13 2.50 ;
        RECT  9.01 3.46 10.05 3.78 ;
        POLYGON  9.69 4.54 8.30 4.54 7.66 3.90 5.72 3.90 5.72 1.86 6.04 1.86
                 6.04 3.58 7.80 3.58 8.44 4.22 9.69 4.22 ;
        RECT  8.60 1.22 9.60 1.54 ;
        POLYGON  8.63 3.63 8.31 3.63 8.31 3.26 6.38 3.26 6.38 2.94 7.90 2.94
                 7.90 1.22 8.22 1.22 8.22 2.94 8.63 2.94 ;
        RECT  4.34 1.22 7.52 1.54 ;
        RECT  4.34 4.22 7.52 4.54 ;
        POLYGON  5.36 2.18 1.56 2.18 1.56 1.22 1.88 1.22 1.88 1.86 5.36 1.86 ;
        RECT  2.96 3.58 5.36 3.90 ;
        RECT  2.96 1.22 3.96 1.54 ;
        RECT  1.56 4.22 3.96 4.54 ;
        POLYGON  2.74 2.98 2.40 2.98 2.40 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 1.86 0.50 1.86 0.50 3.58 2.08 3.58 2.08 2.66 2.74 2.66 ;
    END
END sdffnq_2

MACRO sdffnq_1
    CLASS CORE ;
    FOREIGN sdffnq_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 20.48 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  13.63 3.46 12.64 3.46 12.64 3.68 12.32 3.68 12.32 3.14
                 13.63 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.68 2.66 4.32 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.32 3.04 20.11 3.04 20.11 4.54 19.79 4.54 19.79 3.04
                 19.55 3.04 19.55 1.22 19.87 1.22 19.87 2.72 20.32 2.72 ;
        END
    END q
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.66 5.28 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.66 1.76 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 0.90 19.17 0.90 19.17 1.54 18.85 1.54 18.85 0.90
                 17.79 0.90 17.79 1.14 17.47 1.14 17.47 0.90 10.30 0.90
                 10.30 1.48 9.98 1.48 9.98 0.90 2.58 0.90 2.58 1.54 2.26 1.54
                 2.26 0.90 1.20 0.90 1.20 1.86 0.88 1.86 0.88 0.90 0.00 0.90
                 0.00 -0.90 20.48 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 10.54 4.86 10.54 3.74 10.86 3.74 10.86 4.86
                 17.53 4.86 17.53 3.96 17.85 3.96 17.85 4.86 19.09 4.86
                 19.09 4.22 19.41 4.22 19.41 4.86 20.48 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  18.73 4.54 18.17 4.54 18.17 3.18 17.19 3.18 17.19 2.86
                 18.17 2.86 18.17 1.22 18.49 1.22 18.49 4.22 18.73 4.22 ;
        POLYGON  17.85 2.47 17.53 2.47 17.53 2.28 15.63 2.28 15.63 4.54
                 15.31 4.54 15.31 2.28 14.87 1.84 14.87 1.22 15.19 1.22
                 15.19 1.70 15.45 1.96 17.85 1.96 ;
        RECT  16.09 3.96 17.09 4.28 ;
        RECT  15.69 1.22 16.99 1.54 ;
        RECT  11.97 4.22 14.93 4.54 ;
        POLYGON  14.77 3.90 13.93 3.90 13.93 3.58 14.45 3.58 14.45 2.34
                 14.29 2.18 11.26 2.18 11.26 1.86 14.43 1.86 14.77 2.20 ;
        RECT  11.73 1.22 14.37 1.54 ;
        POLYGON  14.13 2.86 13.81 2.86 13.81 2.82 11.69 2.82 11.69 3.90
                 11.37 3.90 11.37 2.82 9.27 2.82 9.27 3.13 8.95 3.13 8.95 2.50
                 10.62 2.50 10.62 1.22 11.00 1.22 11.00 1.54 10.94 1.54
                 10.94 2.50 14.13 2.50 ;
        RECT  9.01 3.46 10.05 3.78 ;
        POLYGON  9.69 4.54 8.30 4.54 7.66 3.90 5.72 3.90 5.72 1.86 6.04 1.86
                 6.04 3.58 7.80 3.58 8.44 4.22 9.69 4.22 ;
        RECT  8.60 1.22 9.60 1.54 ;
        POLYGON  8.63 3.63 8.31 3.63 8.31 3.26 6.38 3.26 6.38 2.94 7.90 2.94
                 7.90 1.22 8.22 1.22 8.22 2.94 8.63 2.94 ;
        RECT  4.34 1.22 7.52 1.54 ;
        RECT  4.34 4.22 7.52 4.54 ;
        POLYGON  5.36 2.18 1.56 2.18 1.56 1.22 1.88 1.22 1.88 1.86 5.36 1.86 ;
        RECT  2.96 3.58 5.36 3.90 ;
        RECT  2.96 1.22 3.96 1.54 ;
        RECT  1.56 4.22 3.96 4.54 ;
        POLYGON  2.74 2.98 2.40 2.98 2.40 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 1.86 0.50 1.86 0.50 3.58 2.08 3.58 2.08 2.66 2.74 2.66 ;
    END
END sdffnq_1

MACRO sdffn_4
    CLASS CORE ;
    FOREIGN sdffn_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  13.63 3.46 12.64 3.46 12.64 3.68 12.32 3.68 12.32 3.14
                 13.63 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.68 2.66 4.32 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  21.10 3.25 19.33 3.25 19.33 2.93 20.64 2.93 20.64 2.71
                 20.78 2.71 20.78 1.96 18.85 1.96 18.85 1.64 21.10 1.64 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  23.52 4.53 21.42 4.53 21.42 4.21 23.20 4.21 23.20 1.90
                 21.42 1.90 21.42 1.58 23.52 1.58 ;
        END
    END qb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.66 5.28 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.66 1.76 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  23.68 0.90 22.44 0.90 22.44 1.23 22.12 1.23 22.12 0.90
                 19.87 0.90 19.87 1.23 19.55 1.23 19.55 0.90 17.79 0.90
                 17.79 1.14 17.47 1.14 17.47 0.90 10.30 0.90 10.30 1.48
                 9.98 1.48 9.98 0.90 2.58 0.90 2.58 1.54 2.26 1.54 2.26 0.90
                 1.20 0.90 1.20 1.86 0.88 1.86 0.88 0.90 0.00 0.90 0.00 -0.90
                 23.68 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  23.68 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 10.54 4.86 10.54 3.74 10.86 3.74 10.86 4.86
                 17.53 4.86 17.53 3.96 17.85 3.96 17.85 4.86 19.97 4.86
                 19.97 4.79 20.39 4.79 20.39 4.86 23.68 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  22.44 3.89 20.18 3.89 20.18 4.24 18.17 4.24 18.17 3.18
                 17.19 3.18 17.19 2.86 18.17 2.86 18.17 1.22 18.49 1.22
                 18.49 3.92 19.86 3.92 19.86 3.57 22.12 3.57 22.12 2.33
                 22.44 2.33 ;
        POLYGON  17.85 2.47 17.53 2.47 17.53 2.28 15.63 2.28 15.63 4.54
                 15.31 4.54 15.31 2.28 14.87 1.84 14.87 1.22 15.19 1.22
                 15.19 1.70 15.45 1.96 17.85 1.96 ;
        RECT  16.09 3.96 17.09 4.28 ;
        RECT  15.69 1.22 16.99 1.54 ;
        RECT  11.97 4.22 14.93 4.54 ;
        POLYGON  14.77 3.90 13.93 3.90 13.93 3.58 14.45 3.58 14.45 2.34
                 14.29 2.18 11.26 2.18 11.26 1.86 14.43 1.86 14.77 2.20 ;
        RECT  11.73 1.22 14.37 1.54 ;
        POLYGON  14.13 2.86 13.81 2.86 13.81 2.82 11.69 2.82 11.69 3.90
                 11.37 3.90 11.37 2.82 9.27 2.82 9.27 3.13 8.95 3.13 8.95 2.50
                 10.62 2.50 10.62 1.22 11.00 1.22 11.00 1.54 10.94 1.54
                 10.94 2.50 14.13 2.50 ;
        RECT  9.01 3.46 10.05 3.78 ;
        POLYGON  9.69 4.54 8.30 4.54 7.66 3.90 5.72 3.90 5.72 1.86 6.04 1.86
                 6.04 3.58 7.80 3.58 8.44 4.22 9.69 4.22 ;
        RECT  8.60 1.22 9.60 1.54 ;
        POLYGON  8.63 3.63 8.31 3.63 8.31 3.26 6.38 3.26 6.38 2.94 7.90 2.94
                 7.90 1.22 8.22 1.22 8.22 2.94 8.63 2.94 ;
        RECT  4.34 1.22 7.52 1.54 ;
        RECT  4.34 4.22 7.52 4.54 ;
        POLYGON  5.36 2.18 1.56 2.18 1.56 1.22 1.88 1.22 1.88 1.86 5.36 1.86 ;
        RECT  2.96 3.58 5.36 3.90 ;
        RECT  2.96 1.22 3.96 1.54 ;
        RECT  1.56 4.22 3.96 4.54 ;
        POLYGON  2.74 2.98 2.40 2.98 2.40 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 1.86 0.50 1.86 0.50 3.58 2.08 3.58 2.08 2.66 2.74 2.66 ;
    END
END sdffn_4

MACRO sdffn_2
    CLASS CORE ;
    FOREIGN sdffn_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  13.63 3.46 12.64 3.46 12.64 3.68 12.32 3.68 12.32 3.14
                 13.63 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.68 2.66 4.32 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.84  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  19.68 3.04 19.41 3.04 19.41 3.75 19.09 3.75 19.09 3.04
                 18.85 3.04 18.85 1.64 19.17 1.64 19.17 2.72 19.68 2.72 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.96 4.54 20.58 4.54 20.58 4.22 20.64 4.22 20.64 1.64
                 20.25 1.64 20.25 1.32 20.96 1.32 ;
        END
    END qb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.66 5.28 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.66 1.76 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 0.90 19.87 0.90 19.87 1.24 19.55 1.24 19.55 0.90
                 17.79 0.90 17.79 1.14 17.47 1.14 17.47 0.90 10.30 0.90
                 10.30 1.48 9.98 1.48 9.98 0.90 2.58 0.90 2.58 1.54 2.26 1.54
                 2.26 0.90 1.20 0.90 1.20 1.86 0.88 1.86 0.88 0.90 0.00 0.90
                 0.00 -0.90 21.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 10.54 4.86 10.54 3.74 10.86 3.74 10.86 4.86
                 17.53 4.86 17.53 3.96 17.85 3.96 17.85 4.86 21.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.32 3.92 20.18 3.92 20.18 4.54 18.17 4.54 18.17 3.18
                 17.19 3.18 17.19 2.86 18.17 2.86 18.17 1.22 18.49 1.22
                 18.49 4.22 19.86 4.22 19.86 3.60 20.00 3.60 20.00 2.14
                 20.32 2.14 ;
        POLYGON  17.85 2.47 17.53 2.47 17.53 2.28 15.63 2.28 15.63 4.54
                 15.31 4.54 15.31 2.28 14.87 1.84 14.87 1.22 15.19 1.22
                 15.19 1.70 15.45 1.96 17.85 1.96 ;
        RECT  16.09 3.96 17.09 4.28 ;
        RECT  15.69 1.22 16.99 1.54 ;
        RECT  11.97 4.22 14.93 4.54 ;
        POLYGON  14.77 3.90 13.93 3.90 13.93 3.58 14.45 3.58 14.45 2.34
                 14.29 2.18 11.26 2.18 11.26 1.86 14.43 1.86 14.77 2.20 ;
        RECT  11.73 1.22 14.37 1.54 ;
        POLYGON  14.13 2.86 13.81 2.86 13.81 2.82 11.69 2.82 11.69 3.90
                 11.37 3.90 11.37 2.82 9.27 2.82 9.27 3.13 8.95 3.13 8.95 2.50
                 10.62 2.50 10.62 1.22 11.00 1.22 11.00 1.54 10.94 1.54
                 10.94 2.50 14.13 2.50 ;
        RECT  9.01 3.46 10.05 3.78 ;
        POLYGON  9.69 4.54 8.30 4.54 7.66 3.90 5.72 3.90 5.72 1.86 6.04 1.86
                 6.04 3.58 7.80 3.58 8.44 4.22 9.69 4.22 ;
        RECT  8.60 1.22 9.60 1.54 ;
        POLYGON  8.63 3.63 8.31 3.63 8.31 3.26 6.38 3.26 6.38 2.94 7.90 2.94
                 7.90 1.22 8.22 1.22 8.22 2.94 8.63 2.94 ;
        RECT  4.34 1.22 7.52 1.54 ;
        RECT  4.34 4.22 7.52 4.54 ;
        POLYGON  5.36 2.18 1.56 2.18 1.56 1.22 1.88 1.22 1.88 1.86 5.36 1.86 ;
        RECT  2.96 3.58 5.36 3.90 ;
        RECT  2.96 1.22 3.96 1.54 ;
        RECT  1.56 4.22 3.96 4.54 ;
        POLYGON  2.74 2.98 2.40 2.98 2.40 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 1.86 0.50 1.86 0.50 3.58 2.08 3.58 2.08 2.66 2.74 2.66 ;
    END
END sdffn_2

MACRO sdffn_1
    CLASS CORE ;
    FOREIGN sdffn_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  13.63 3.46 12.64 3.46 12.64 3.68 12.32 3.68 12.32 3.14
                 13.63 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.68 2.66 4.32 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.35  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  19.68 3.04 19.41 3.04 19.41 3.90 19.09 3.90 19.09 3.04
                 18.85 3.04 18.85 1.22 19.17 1.22 19.17 2.72 19.68 2.72 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.21  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.96 4.54 20.58 4.54 20.58 4.22 20.64 4.22 20.64 1.54
                 20.25 1.54 20.25 1.22 20.96 1.22 ;
        END
    END qb
    PIN sdi
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.66 5.28 3.04 ;
        END
    END sdi
    PIN se
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.66 1.76 3.04 ;
        END
    END se
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 0.90 19.87 0.90 19.87 1.54 19.55 1.54 19.55 0.90
                 17.79 0.90 17.79 1.54 17.47 1.54 17.47 0.90 10.30 0.90
                 10.30 1.48 9.98 1.48 9.98 0.90 2.58 0.90 2.58 1.54 2.26 1.54
                 2.26 0.90 1.20 0.90 1.20 1.86 0.88 1.86 0.88 0.90 0.00 0.90
                 0.00 -0.90 21.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 10.54 4.86 10.54 3.74 10.86 3.74 10.86 4.86
                 17.53 4.86 17.53 3.96 17.85 3.96 17.85 4.86 21.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.32 3.77 20.18 3.77 20.18 4.54 18.17 4.54 18.17 3.18
                 17.19 3.18 17.19 2.86 18.17 2.86 18.17 1.22 18.49 1.22
                 18.49 4.22 19.86 4.22 19.86 3.45 20.00 3.45 20.00 2.14
                 20.32 2.14 ;
        POLYGON  17.85 2.47 17.53 2.47 17.53 2.28 15.63 2.28 15.63 4.54
                 15.31 4.54 15.31 2.28 14.87 1.84 14.87 1.22 15.19 1.22
                 15.19 1.70 15.45 1.96 17.85 1.96 ;
        RECT  16.09 3.96 17.09 4.28 ;
        RECT  15.69 1.22 16.99 1.54 ;
        RECT  11.97 4.22 14.93 4.54 ;
        POLYGON  14.77 3.90 13.93 3.90 13.93 3.58 14.45 3.58 14.45 2.34
                 14.29 2.18 11.26 2.18 11.26 1.86 14.43 1.86 14.77 2.20 ;
        RECT  11.73 1.22 14.37 1.54 ;
        POLYGON  14.13 2.86 13.81 2.86 13.81 2.82 11.69 2.82 11.69 3.90
                 11.37 3.90 11.37 2.82 9.27 2.82 9.27 3.13 8.95 3.13 8.95 2.50
                 10.62 2.50 10.62 1.22 11.00 1.22 11.00 1.54 10.94 1.54
                 10.94 2.50 14.13 2.50 ;
        RECT  9.01 3.46 10.05 3.78 ;
        POLYGON  9.69 4.54 8.30 4.54 7.66 3.90 5.72 3.90 5.72 1.86 6.04 1.86
                 6.04 3.58 7.80 3.58 8.44 4.22 9.69 4.22 ;
        RECT  8.60 1.22 9.60 1.54 ;
        POLYGON  8.63 3.63 8.31 3.63 8.31 3.26 6.38 3.26 6.38 2.94 7.90 2.94
                 7.90 1.22 8.22 1.22 8.22 2.94 8.63 2.94 ;
        RECT  4.34 1.22 7.52 1.54 ;
        RECT  4.34 4.22 7.52 4.54 ;
        POLYGON  5.36 2.18 1.56 2.18 1.56 1.22 1.88 1.22 1.88 1.86 5.36 1.86 ;
        RECT  2.96 3.58 5.36 3.90 ;
        RECT  2.96 1.22 3.96 1.54 ;
        RECT  1.56 4.22 3.96 4.54 ;
        POLYGON  2.74 2.98 2.40 2.98 2.40 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 1.86 0.50 1.86 0.50 3.58 2.08 3.58 2.08 2.66 2.74 2.66 ;
    END
END sdffn_1

MACRO or4_8
    CLASS CORE ;
    FOREIGN or4_8 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.72 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.32  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 1.76 0.48 2.40 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.32  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.08 3.04 2.72 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.32  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 1.86 6.88 2.50 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.32  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.08 4.22 2.40 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.91  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.08 4.54 7.82 4.54 7.82 4.22 11.68 4.22 11.68 4.00
                 11.92 4.00 11.92 2.18 7.82 2.18 7.82 1.22 8.14 1.22 8.14 1.86
                 12.24 1.86 12.24 4.22 14.08 4.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  14.72 0.90 7.46 0.90 7.46 1.54 7.14 1.54 7.14 0.90 4.32 0.90
                 4.32 1.54 4.00 1.54 4.00 0.90 3.64 0.90 3.64 1.54 3.32 1.54
                 3.32 0.90 0.00 0.90 0.00 -0.90 14.72 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  14.72 6.66 0.00 6.66 0.00 4.86 3.66 4.86 3.66 4.22 3.98 4.22
                 3.98 4.86 14.72 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  8.52 1.22 14.42 1.54 ;
        POLYGON  11.60 3.26 11.28 3.26 11.28 2.94 9.98 2.94 9.98 3.26 5.74 3.26
                 5.74 1.54 4.70 1.54 4.70 1.22 6.76 1.22 6.76 1.54 6.06 1.54
                 6.06 2.94 9.66 2.94 9.66 2.62 11.60 2.62 ;
        POLYGON  10.62 3.90 1.58 3.90 1.58 3.26 0.50 3.26 0.50 4.54 0.18 4.54
                 0.18 2.94 0.80 2.94 0.80 1.22 2.94 1.22 2.94 1.54 1.12 1.54
                 1.12 2.94 1.90 2.94 1.90 3.58 10.30 3.58 10.30 3.26 10.62 3.26 ;
        RECT  4.36 4.22 6.76 4.54 ;
        RECT  0.88 4.22 3.28 4.54 ;
    END
END or4_8

MACRO or4_4
    CLASS CORE ;
    FOREIGN or4_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.24 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 1.76 0.48 2.40 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 1.76 2.72 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 1.79 4.32 2.43 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.08 2.82 2.40 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.19  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.86 4.54 5.74 4.54 5.74 4.22 7.84 4.22 7.84 4.00 8.10 4.00
                 8.10 2.18 5.31 2.18 5.31 1.86 8.42 1.86 8.42 4.22 8.86 4.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  10.24 0.90 9.81 0.90 9.81 1.54 9.49 1.54 9.49 0.90 4.23 0.90
                 4.23 1.19 3.91 1.19 3.91 0.90 2.83 0.90 2.83 1.19 2.51 1.19
                 2.51 0.90 2.15 0.90 2.15 1.18 1.83 1.18 1.83 0.90 0.00 0.90
                 0.00 -0.90 10.24 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  10.24 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.26 2.58 4.26
                 2.58 4.86 5.04 4.86 5.04 4.22 5.36 4.22 5.36 4.86 9.24 4.86
                 9.24 4.22 9.56 4.22 9.56 4.86 10.24 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  4.61 1.22 9.11 1.54 ;
        POLYGON  7.78 3.26 7.46 3.26 7.46 2.94 6.50 2.94 6.50 3.26 3.14 3.26
                 3.14 1.44 3.21 1.44 3.21 1.22 3.53 1.22 3.53 1.76 3.46 1.76
                 3.46 2.94 6.18 2.94 6.18 2.62 7.78 2.62 ;
        POLYGON  7.14 3.90 0.50 3.90 0.50 4.54 0.18 4.54 0.18 3.58 0.80 3.58
                 0.80 1.22 1.45 1.22 1.45 1.54 1.12 1.54 1.12 3.58 6.82 3.58
                 6.82 3.26 7.14 3.26 ;
        RECT  2.96 4.22 3.96 4.54 ;
        RECT  0.88 4.22 1.88 4.54 ;
    END
END or4_4

MACRO or4_2
    CLASS CORE ;
    FOREIGN or4_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.96 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 1.76 0.48 2.40 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 1.76 2.72 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 1.79 4.32 2.43 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.08 2.82 2.40 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.16  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.14 4.54 5.02 4.54 5.02 4.22 7.20 4.22 7.20 4.00 7.38 4.00
                 7.38 2.18 5.38 2.18 5.38 1.86 7.70 1.86 7.70 4.22 8.14 4.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.96 0.90 4.32 0.90 4.32 1.18 4.00 1.18 4.00 0.90 2.92 0.90
                 2.92 1.19 2.60 1.19 2.60 0.90 2.24 0.90 2.24 1.18 1.92 1.18
                 1.92 0.90 0.00 0.90 0.00 -0.90 8.96 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  8.96 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.22 2.58 4.22
                 2.58 4.86 8.96 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  4.68 1.22 8.48 1.54 ;
        POLYGON  7.06 3.26 6.74 3.26 6.74 2.94 5.78 2.94 5.78 3.26 3.14 3.26
                 3.14 1.44 3.30 1.44 3.30 1.22 3.62 1.22 3.62 1.76 3.46 1.76
                 3.46 2.94 5.46 2.94 5.46 2.62 7.06 2.62 ;
        POLYGON  6.42 3.90 0.50 3.90 0.50 4.54 0.18 4.54 0.18 3.58 0.80 3.58
                 0.80 1.22 1.54 1.22 1.54 1.54 1.12 1.54 1.12 3.58 6.10 3.58
                 6.10 3.26 6.42 3.26 ;
        RECT  2.96 4.22 3.96 4.54 ;
        RECT  0.88 4.22 1.88 4.54 ;
    END
END or4_2

MACRO or4_1
    CLASS CORE ;
    FOREIGN or4_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.04 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.08 0.48 2.72 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 1.76 2.72 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 1.86 4.32 2.50 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.08 2.82 2.40 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  6.88 4.54 5.02 4.54 5.02 4.22 6.56 4.22 6.56 2.18 5.14 2.18
                 5.14 1.86 6.88 1.86 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 7.04 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.04 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.22 2.58 4.22
                 2.58 4.86 7.04 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  4.44 1.22 6.84 1.54 ;
        POLYGON  6.24 2.94 5.08 2.94 5.08 3.26 3.14 3.26 3.14 1.54 2.26 1.54
                 2.26 1.22 3.98 1.22 3.98 1.54 3.46 1.54 3.46 2.94 4.76 2.94
                 4.76 2.62 6.24 2.62 ;
        POLYGON  5.72 3.90 0.50 3.90 0.50 4.54 0.18 4.54 0.18 3.58 0.80 3.58
                 0.80 1.54 0.18 1.54 0.18 1.22 1.90 1.22 1.90 1.54 1.12 1.54
                 1.12 3.58 5.40 3.58 5.40 3.26 5.72 3.26 ;
        RECT  2.96 4.22 3.96 4.54 ;
        RECT  0.88 4.22 1.88 4.54 ;
    END
END or4_1

MACRO or3_8
    CLASS CORE ;
    FOREIGN or3_8 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 1.90 0.90 2.54 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 1.90 2.40 2.54 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 1.98 3.68 2.62 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.93  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  6.54 4.54 6.22 4.54 6.22 2.40 4.96 2.40 4.96 3.90 4.90 3.90
                 4.90 4.54 4.58 4.54 4.58 3.58 4.64 3.58 4.64 1.54 4.58 1.54
                 4.58 1.22 4.96 1.22 4.96 2.08 6.22 2.08 6.22 1.33 6.54 1.33 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 0.90 7.24 0.90 7.24 1.66 6.92 1.66 6.92 0.90 5.60 0.90
                 5.60 1.66 5.28 1.66 5.28 0.90 3.89 0.90 3.89 1.54 3.57 1.54
                 3.57 0.90 2.22 0.90 2.22 1.54 1.90 1.54 1.90 0.90 0.84 0.90
                 0.84 1.54 0.52 1.54 0.52 0.90 0.00 0.90 0.00 -0.90 7.68 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 6.66 0.00 6.66 0.00 4.86 3.75 4.86 3.75 3.58 4.07 3.58
                 4.07 4.86 5.28 4.86 5.28 3.58 5.60 3.58 5.60 4.86 6.92 4.86
                 6.92 3.58 7.24 3.58 7.24 4.86 7.68 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.32 3.26 0.50 3.26 0.50 4.54 0.18 4.54 0.18 2.94 1.22 2.94
                 1.22 1.22 1.54 1.22 1.54 2.94 2.72 2.94 2.72 1.54 2.60 1.54
                 2.60 1.22 3.04 1.22 3.04 2.94 4.00 2.94 4.00 2.13 4.32 2.13 ;
        RECT  2.26 3.58 3.26 4.54 ;
        RECT  0.88 3.58 1.88 4.54 ;
    END
END or3_8

MACRO or3_4
    CLASS CORE ;
    FOREIGN or3_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 1.90 0.90 2.54 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 1.90 2.40 2.54 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 1.98 3.68 2.62 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.97  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.96 3.90 4.90 3.90 4.90 4.54 4.58 4.54 4.58 3.58 4.64 3.58
                 4.64 1.54 4.58 1.54 4.58 1.22 4.96 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 0.90 5.60 0.90 5.60 1.66 5.28 1.66 5.28 0.90 3.89 0.90
                 3.89 1.54 3.57 1.54 3.57 0.90 2.22 0.90 2.22 1.54 1.90 1.54
                 1.90 0.90 0.84 0.90 0.84 1.54 0.52 1.54 0.52 0.90 0.00 0.90
                 0.00 -0.90 6.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 6.66 0.00 6.66 0.00 4.86 3.75 4.86 3.75 3.58 4.07 3.58
                 4.07 4.86 5.28 4.86 5.28 3.58 5.60 3.58 5.60 4.86 6.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.32 3.26 0.50 3.26 0.50 4.54 0.18 4.54 0.18 2.94 1.22 2.94
                 1.22 1.22 1.54 1.22 1.54 2.94 2.72 2.94 2.72 1.54 2.60 1.54
                 2.60 1.22 3.04 1.22 3.04 2.94 4.00 2.94 4.00 2.13 4.32 2.13 ;
        RECT  2.26 3.58 3.26 4.54 ;
        RECT  0.88 3.58 1.88 4.54 ;
    END
END or3_4

MACRO or3_2
    CLASS CORE ;
    FOREIGN or3_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 1.90 0.80 2.54 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 1.90 2.40 2.54 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.24 2.08 3.68 2.61 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.96 4.54 4.62 4.54 4.62 4.22 4.64 4.22 4.64 1.54 4.14 1.54
                 4.14 1.22 4.96 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 0.90 3.60 0.90 3.60 1.54 3.28 1.54 3.28 0.90 0.74 0.90
                 0.74 1.54 0.42 1.54 0.42 0.90 0.00 0.90 0.00 -0.90 5.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 6.66 0.00 6.66 0.00 4.86 3.76 4.86 3.76 4.22 4.08 4.22
                 4.08 4.86 5.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.32 3.25 0.50 3.25 0.50 4.54 0.18 4.54 0.18 2.93 1.12 2.93
                 1.12 1.22 2.83 1.22 2.83 1.54 1.44 1.54 1.44 2.93 4.00 2.93
                 4.00 2.12 4.32 2.12 ;
        RECT  2.26 3.58 3.26 4.54 ;
        RECT  0.88 3.58 1.88 4.54 ;
    END
END or3_2

MACRO or3_1
    CLASS CORE ;
    FOREIGN or3_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 1.90 0.90 2.40 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 1.90 2.40 2.54 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 1.90 3.68 2.54 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.96 4.54 4.58 4.54 4.58 4.22 4.64 4.22 4.64 1.54 4.58 1.54
                 4.58 1.22 4.96 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 0.90 3.89 0.90 3.89 1.54 3.57 1.54 3.57 0.90 2.22 0.90
                 2.22 1.54 1.90 1.54 1.90 0.90 0.84 0.90 0.84 1.54 0.52 1.54
                 0.52 0.90 0.00 0.90 0.00 -0.90 5.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 6.66 0.00 6.66 0.00 4.86 3.75 4.86 3.75 4.28 4.07 4.28
                 4.07 4.86 5.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.32 3.25 0.50 3.25 0.50 4.54 0.18 4.54 0.18 2.93 1.22 2.93
                 1.22 1.22 1.54 1.22 1.54 2.93 2.72 2.93 2.72 1.54 2.60 1.54
                 2.60 1.22 3.04 1.22 3.04 2.93 4.00 2.93 4.00 2.11 4.32 2.11 ;
        RECT  2.26 3.58 3.26 4.54 ;
        RECT  0.88 3.58 1.88 4.54 ;
    END
END or3_1

MACRO or2a_8
    CLASS CORE ;
    FOREIGN or2a_8 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.60 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.45  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.72 1.12 3.36 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.32  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 1.86 4.96 2.50 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.93  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.94 4.54 7.62 4.54 7.62 2.40 6.30 2.40 6.30 4.54 5.98 4.54
                 5.98 2.40 5.92 2.40 5.92 2.08 5.98 2.08 5.98 1.22 6.30 1.22
                 6.30 2.08 7.62 2.08 7.62 1.22 7.94 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  9.60 0.90 8.64 0.90 8.64 1.54 8.32 1.54 8.32 0.90 7.11 0.90
                 7.11 1.54 6.79 1.54 6.79 0.90 5.44 0.90 5.44 1.54 5.12 1.54
                 5.12 0.90 1.20 0.90 1.20 1.54 0.88 1.54 0.88 0.90 0.00 0.90
                 0.00 -0.90 9.60 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  9.60 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.26 1.20 4.26
                 1.20 4.86 5.16 4.86 5.16 3.57 5.48 3.57 5.48 4.86 6.80 4.86
                 6.80 3.57 7.12 3.57 7.12 4.86 8.32 4.86 8.32 3.56 8.64 3.56
                 8.64 4.86 9.60 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  5.60 3.25 3.28 3.25 3.28 3.89 2.96 3.89 2.96 3.25 1.88 3.25
                 1.88 4.54 1.56 4.54 1.56 2.93 2.96 2.93 2.96 1.54 1.56 1.54
                 1.56 1.22 4.66 1.22 4.66 1.54 3.28 1.54 3.28 2.93 5.28 2.93
                 5.28 2.12 5.60 2.12 ;
        POLYGON  4.66 4.54 2.26 4.54 2.26 3.57 2.58 3.57 2.58 4.22 4.34 4.22
                 4.34 3.57 4.66 3.57 ;
        POLYGON  2.28 2.22 0.48 2.22 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 1.90 2.28 1.90 ;
    END
END or2a_8

MACRO or2a_4
    CLASS CORE ;
    FOREIGN or2a_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.45  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.72 1.12 3.36 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.24 1.86 3.68 2.50 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.02  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 1.22 4.96 4.54 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 0.90 3.78 0.90 3.78 1.54 3.46 1.54 3.46 0.90 2.22 0.90
                 2.22 1.54 1.90 1.54 1.90 0.90 1.20 0.90 1.20 1.54 0.88 1.54
                 0.88 0.90 0.00 0.90 0.00 -0.90 6.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.26 1.20 4.26
                 1.20 4.86 3.75 4.86 3.75 4.22 4.07 4.22 4.07 4.86 6.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.32 3.25 1.88 3.25 1.88 4.54 1.56 4.54 1.56 2.93 2.60 2.93
                 2.60 1.22 2.92 1.22 2.92 2.93 4.00 2.93 4.00 2.12 4.32 2.12 ;
        RECT  2.26 3.58 3.26 4.54 ;
        POLYGON  2.28 2.22 0.48 2.22 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 1.90 2.28 1.90 ;
    END
END or2a_4

MACRO or2a_2
    CLASS CORE ;
    FOREIGN or2a_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.45  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.72 1.12 3.36 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.24 1.86 3.68 2.50 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.96 4.13 4.90 4.13 4.90 4.54 4.58 4.54 4.58 3.81 4.64 3.81
                 4.64 1.54 4.58 1.54 4.58 1.22 4.96 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 0.90 3.78 0.90 3.78 1.54 3.46 1.54 3.46 0.90 2.22 0.90
                 2.22 1.54 1.90 1.54 1.90 0.90 1.20 0.90 1.20 1.54 0.88 1.54
                 0.88 0.90 0.00 0.90 0.00 -0.90 5.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.26 1.20 4.26
                 1.20 4.86 3.75 4.86 3.75 4.22 4.07 4.22 4.07 4.86 5.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.32 3.25 1.88 3.25 1.88 4.54 1.56 4.54 1.56 2.93 2.60 2.93
                 2.60 1.22 2.92 1.22 2.92 2.93 4.00 2.93 4.00 2.12 4.32 2.12 ;
        RECT  2.26 3.58 3.26 4.54 ;
        POLYGON  2.28 2.22 0.48 2.22 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 1.90 2.28 1.90 ;
    END
END or2a_2

MACRO or2a_1
    CLASS CORE ;
    FOREIGN or2a_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.45  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.72 1.12 3.36 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 1.86 3.68 2.50 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.96 4.54 4.58 4.54 4.58 4.22 4.64 4.22 4.64 1.54 4.58 1.54
                 4.58 1.22 4.96 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 0.90 3.91 0.90 3.91 1.54 3.59 1.54 3.59 0.90 2.22 0.90
                 2.22 1.54 1.90 1.54 1.90 0.90 1.20 0.90 1.20 1.54 0.88 1.54
                 0.88 0.90 0.00 0.90 0.00 -0.90 5.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.26 1.20 4.26
                 1.20 4.86 3.75 4.86 3.75 4.27 4.07 4.27 4.07 4.86 5.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.32 3.25 1.88 3.25 1.88 4.54 1.56 4.54 1.56 2.93 2.60 2.93
                 2.60 1.22 2.92 1.22 2.92 2.93 4.00 2.93 4.00 2.12 4.32 2.12 ;
        RECT  2.26 3.58 3.26 4.54 ;
        POLYGON  2.28 2.22 0.48 2.22 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 1.90 2.28 1.90 ;
    END
END or2a_1

MACRO or2_8
    CLASS CORE ;
    FOREIGN or2_8 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.32 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.32  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.90 1.12 2.54 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.32  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 1.86 3.04 2.50 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.99  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  6.41 4.54 6.09 4.54 6.09 2.40 4.92 2.40 4.92 4.54 4.60 4.54
                 4.60 1.22 4.92 1.22 4.92 2.08 6.09 2.08 6.09 1.22 6.41 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 0.90 7.30 0.90 7.30 1.54 6.98 1.54 6.98 0.90 5.62 0.90
                 5.62 1.54 5.30 1.54 5.30 0.90 4.06 0.90 4.06 1.54 3.74 1.54
                 3.74 0.90 0.00 0.90 0.00 -0.90 8.32 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 6.66 0.00 6.66 0.00 4.86 3.78 4.86 3.78 3.57 4.10 3.57
                 4.10 4.86 5.30 4.86 5.30 3.57 5.62 3.57 5.62 4.86 6.98 4.86
                 6.98 4.22 7.30 4.22 7.30 4.86 8.32 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.22 3.25 1.90 3.25 1.90 3.89 1.58 3.89 1.58 3.25 0.50 3.25
                 0.50 4.54 0.16 4.54 0.16 1.22 3.28 1.22 3.28 1.54 0.48 1.54
                 0.48 2.93 3.90 2.93 3.90 2.12 4.22 2.12 ;
        POLYGON  3.28 4.54 0.88 4.54 0.88 3.57 1.20 3.57 1.20 4.22 2.96 4.22
                 2.96 3.57 3.28 3.57 ;
    END
END or2_8

MACRO or2_4
    CLASS CORE ;
    FOREIGN or2_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 1.90 0.48 2.54 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.85 1.86 2.40 2.40 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.97  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.68 4.54 3.20 4.54 3.20 4.22 3.36 4.22 3.36 1.54 3.20 1.54
                 3.20 1.22 3.68 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 0.90 2.36 0.90 2.36 1.54 2.04 1.54 2.04 0.90 0.84 0.90
                 0.84 1.19 0.52 1.19 0.52 0.90 0.00 0.90 0.00 -0.90 5.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 6.66 0.00 6.66 0.00 4.86 2.44 4.86 2.44 4.22 2.76 4.22
                 2.76 4.86 5.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  3.04 3.24 0.50 3.24 0.50 4.54 0.18 4.54 0.18 2.92 1.21 2.92
                 1.21 1.22 1.54 1.22 1.54 1.54 1.53 1.54 1.53 2.92 2.72 2.92
                 2.72 2.12 3.04 2.12 ;
        RECT  0.88 3.57 1.88 4.54 ;
    END
END or2_4

MACRO or2_2
    CLASS CORE ;
    FOREIGN or2_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.84 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 1.90 0.48 2.54 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.85 1.86 2.40 2.41 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.68 4.54 3.20 4.54 3.20 4.22 3.36 4.22 3.36 1.54 3.20 1.54
                 3.20 1.22 3.68 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  3.84 0.90 2.36 0.90 2.36 1.54 2.04 1.54 2.04 0.90 0.84 0.90
                 0.84 1.19 0.52 1.19 0.52 0.90 0.00 0.90 0.00 -0.90 3.84 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  3.84 6.66 0.00 6.66 0.00 4.86 2.44 4.86 2.44 4.22 2.76 4.22
                 2.76 4.86 3.84 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  3.04 3.24 0.50 3.24 0.50 4.54 0.18 4.54 0.18 2.92 1.21 2.92
                 1.21 1.22 1.54 1.22 1.54 1.54 1.53 1.54 1.53 2.92 2.72 2.92
                 2.72 2.12 3.04 2.12 ;
        RECT  0.88 3.57 1.88 4.54 ;
    END
END or2_2

MACRO or2_1
    CLASS CORE ;
    FOREIGN or2_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.84 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 1.90 0.48 2.54 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 1.86 2.40 2.50 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.68 4.54 3.20 4.54 3.20 4.22 3.36 4.22 3.36 1.54 3.20 1.54
                 3.20 1.22 3.68 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  3.84 0.90 2.82 0.90 2.82 1.54 1.92 1.54 1.92 0.90 0.84 0.90
                 0.84 1.19 0.52 1.19 0.52 0.90 0.00 0.90 0.00 -0.90 3.84 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  3.84 6.66 0.00 6.66 0.00 4.86 2.37 4.86 2.37 4.28 2.69 4.28
                 2.69 4.86 3.84 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  3.04 3.25 0.50 3.25 0.50 4.54 0.18 4.54 0.18 2.93 1.22 2.93
                 1.22 1.22 1.54 1.22 1.54 2.93 2.72 2.93 2.72 2.12 3.04 2.12 ;
        RECT  0.88 3.57 1.88 4.54 ;
    END
END or2_1

MACRO oai33_4
    CLASS CORE ;
    FOREIGN oai33_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.16 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.40 6.88 3.04 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.62 1.12 3.26 ;
        END
    END d
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.40 2.62 10.72 3.26 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  8.48 2.62 8.80 3.26 ;
        END
    END b
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.62 3.04 3.26 ;
        END
    END e
    PIN f
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.62 4.96 3.26 ;
        END
    END f
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.46 3.90 6.06 3.90 6.06 4.54 5.74 4.54 5.74 3.90 4.34 3.90
                 4.34 3.58 5.74 3.58 5.74 2.18 0.18 2.18 0.18 1.22 0.50 1.22
                 0.50 1.86 6.06 1.86 6.06 2.72 6.24 2.72 6.24 3.04 6.06 3.04
                 6.06 3.58 7.46 3.58 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 12.16 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  12.16 6.66 0.00 6.66 0.00 4.86 10.60 4.86 10.60 4.22
                 10.92 4.22 10.92 4.86 12.16 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  0.88 1.22 11.62 1.54 ;
        POLYGON  11.62 4.54 11.30 4.54 11.30 3.90 10.22 3.90 10.22 4.54
                 9.90 4.54 9.90 3.90 8.52 3.90 8.52 3.58 11.62 3.58 ;
        POLYGON  9.54 4.54 6.44 4.54 6.44 4.22 7.82 4.22 7.82 3.58 8.14 3.58
                 8.14 4.22 9.54 4.22 ;
        POLYGON  5.36 4.54 3.66 4.54 3.66 3.90 2.26 3.90 2.26 3.58 3.98 3.58
                 3.98 4.22 5.36 4.22 ;
        POLYGON  3.28 4.54 0.18 4.54 0.18 3.58 0.50 3.58 0.50 4.22 1.58 4.22
                 1.58 3.58 1.90 3.58 1.90 4.22 3.28 4.22 ;
    END
END oai33_4

MACRO oai33_2
    CLASS CORE ;
    FOREIGN oai33_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.40 6.88 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 2.40 5.60 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.40 4.32 3.04 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.62 1.12 3.26 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.62 2.40 3.26 ;
        END
    END e
    PIN f
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.62 3.04 3.26 ;
        END
    END f
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.97  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.96 4.54 3.64 4.54 3.64 3.84 3.36 3.84 3.36 2.18 0.46 2.18
                 0.46 1.22 0.78 1.22 0.78 1.86 3.68 1.86 3.68 3.52 3.96 3.52 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 7.68 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 6.40 4.86 6.40 4.22 6.72 4.22 6.72 4.86 7.68 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  1.16 1.22 7.42 1.54 ;
        POLYGON  7.42 4.54 7.10 4.54 7.10 3.90 6.04 3.90 6.04 4.54 5.72 4.54
                 5.72 3.58 7.42 3.58 ;
        RECT  4.34 3.58 5.34 4.54 ;
        POLYGON  3.26 4.54 2.26 4.54 2.26 3.58 2.58 3.58 2.58 4.22 3.26 4.22 ;
        POLYGON  1.88 4.54 1.56 4.54 1.56 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 3.58 1.88 3.58 ;
    END
END oai33_2

MACRO oai33_1
    CLASS CORE ;
    FOREIGN oai33_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.72 6.88 3.36 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 2.72 5.60 3.36 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.72 4.64 3.04 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.72 1.12 3.36 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.72 2.40 3.36 ;
        END
    END e
    PIN f
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.04 3.36 ;
        END
    END f
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.21  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.96 4.54 3.64 4.54 3.64 3.84 3.36 3.84 3.36 2.40 0.46 2.40
                 0.46 1.22 0.78 1.22 0.78 2.08 2.62 2.08 2.62 1.86 2.94 1.86
                 2.94 2.08 3.68 2.08 3.68 3.52 3.96 3.52 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 7.68 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 7.68 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  1.16 1.22 7.42 1.54 ;
        RECT  5.72 4.22 7.42 4.54 ;
        RECT  4.34 4.22 5.34 4.54 ;
        RECT  2.26 4.22 3.26 4.54 ;
        RECT  0.18 4.22 1.88 4.54 ;
    END
END oai33_1

MACRO oai32_4
    CLASS CORE ;
    FOREIGN oai32_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.24 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  8.48 2.40 8.80 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.62 6.88 3.26 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.62 4.96 3.26 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.62 1.12 3.26 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.62 3.04 3.26 ;
        END
    END e
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.29  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  5.38 3.90 3.98 3.90 3.98 4.54 3.66 4.54 3.66 3.90 2.26 3.90
                 2.26 3.58 3.66 3.58 3.66 2.18 0.48 2.18 0.48 2.40 0.16 2.40
                 0.16 1.86 0.18 1.86 0.18 1.22 0.50 1.22 0.50 1.86 3.98 1.86
                 3.98 3.58 5.38 3.58 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 10.24 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  10.24 6.66 0.00 6.66 0.00 4.86 8.52 4.86 8.52 4.22 8.84 4.22
                 8.84 4.86 10.24 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  0.88 1.22 9.54 1.54 ;
        POLYGON  9.54 4.54 9.22 4.54 9.22 3.90 8.14 3.90 8.14 4.54 7.14 4.54
                 7.14 3.90 5.74 3.90 5.74 3.58 7.46 3.58 7.46 4.22 7.82 4.22
                 7.82 3.58 9.54 3.58 ;
        RECT  4.36 4.22 6.76 4.54 ;
        POLYGON  3.28 4.54 0.18 4.54 0.18 3.58 0.50 3.58 0.50 4.22 1.58 4.22
                 1.58 3.58 1.90 3.58 1.90 4.22 3.28 4.22 ;
    END
END oai32_4

MACRO oai32_2
    CLASS CORE ;
    FOREIGN oai32_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 2.40 5.60 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.94 2.40 4.32 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.62 3.04 3.26 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.62 1.12 3.26 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.62 1.76 3.26 ;
        END
    END e
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.29  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  2.58 4.54 2.26 4.54 2.26 3.86 2.08 3.86 2.08 2.18 1.24 2.18
                 1.24 1.86 2.40 1.86 2.40 3.57 2.58 3.57 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 6.40 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 6.66 0.00 6.66 0.00 4.86 5.02 4.86 5.02 4.22 5.34 4.22
                 5.34 4.86 6.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  0.46 1.22 6.04 1.54 ;
        POLYGON  6.04 4.54 5.72 4.54 5.72 3.90 4.66 3.90 4.66 4.54 4.34 4.54
                 4.34 3.58 6.04 3.58 ;
        POLYGON  3.96 4.54 2.96 4.54 2.96 3.58 3.28 3.58 3.28 4.22 3.64 4.22
                 3.64 3.58 3.96 3.58 ;
        POLYGON  1.88 4.54 0.18 4.54 0.18 3.58 0.50 3.58 0.50 4.22 1.88 4.22 ;
    END
END oai32_2

MACRO oai32_1
    CLASS CORE ;
    FOREIGN oai32_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 2.72 5.60 3.36 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.94 2.72 4.32 3.36 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.04 3.36 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.72 1.12 3.36 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.72 1.76 3.36 ;
        END
    END e
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.72  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  2.58 4.06 2.26 4.06 2.26 3.94 2.08 3.94 2.08 2.40 1.24 2.40
                 1.24 1.86 1.56 1.86 1.56 2.08 2.40 2.08 2.40 3.65 2.58 3.65 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 6.40 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 6.40 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  0.46 1.22 6.04 1.54 ;
        RECT  4.34 4.22 6.04 4.54 ;
        RECT  2.96 4.22 3.96 4.54 ;
        RECT  0.18 4.22 1.88 4.54 ;
    END
END oai32_1

MACRO oai31_4
    CLASS CORE ;
    FOREIGN oai31_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.62 6.88 3.26 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.62 4.96 3.26 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.62 2.40 3.26 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.62 1.12 3.26 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.30 3.90 1.90 3.90 1.90 4.54 1.58 4.54 1.58 3.90 0.50 3.90
                 0.50 4.54 0.16 4.54 0.16 1.86 0.18 1.86 0.18 1.22 0.50 1.22
                 0.50 1.86 1.90 1.86 1.90 2.18 0.48 2.18 0.48 3.58 3.30 3.58 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 7.68 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 6.44 4.86 6.44 4.22 6.76 4.22 6.76 4.86 7.68 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  0.88 1.22 7.46 1.54 ;
        POLYGON  7.46 4.54 7.14 4.54 7.14 3.90 6.06 3.90 6.06 4.54 5.74 4.54
                 5.74 3.90 5.38 3.90 5.38 4.54 5.06 4.54 5.06 3.90 3.66 3.90
                 3.66 3.58 7.46 3.58 ;
        RECT  2.28 4.22 4.68 4.54 ;
    END
END oai31_4

MACRO oai31_2
    CLASS CORE ;
    FOREIGN oai31_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.40 4.32 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.40 3.04 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.40 1.76 3.04 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.40 1.12 3.04 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.84  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.44 4.06 0.16 4.06 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 3.74 1.44 3.74 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 0.90 4.66 0.90 4.66 1.54 4.34 1.54 4.34 0.90 0.00 0.90
                 0.00 -0.90 5.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 6.66 0.00 6.66 0.00 4.86 3.88 4.86 3.88 4.22 4.20 4.22
                 4.20 4.86 5.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.90 4.54 4.58 4.54 4.58 3.90 3.52 3.90 3.52 4.54 3.20 4.54
                 3.20 3.58 4.90 3.58 ;
        RECT  0.88 1.22 3.96 1.54 ;
        RECT  1.82 3.58 2.82 4.54 ;
    END
END oai31_2

MACRO oai31_1
    CLASS CORE ;
    FOREIGN oai31_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.72 4.32 3.36 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.04 3.36 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.72 1.76 3.36 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.72 1.12 3.36 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.32  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.44 4.06 0.16 4.06 0.16 1.34 0.50 1.34 0.50 1.66 0.48 1.66
                 0.48 3.74 1.44 3.74 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 0.90 4.66 0.90 4.66 1.66 4.34 1.66 4.34 0.90 0.00 0.90
                 0.00 -0.90 5.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 5.12 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  3.20 4.22 4.90 4.54 ;
        RECT  0.88 1.22 3.96 1.54 ;
        RECT  1.82 4.22 2.82 4.54 ;
    END
END oai31_1

MACRO oai22_4
    CLASS CORE ;
    FOREIGN oai22_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.40 6.88 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.40 4.96 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.62 1.12 3.26 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.62 3.04 3.04 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.29  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  5.38 3.68 3.98 3.68 3.98 4.54 3.66 4.54 3.66 3.68 2.26 3.68
                 2.26 3.36 3.66 3.36 3.66 2.22 0.18 2.22 0.18 1.22 0.50 1.22
                 0.50 1.90 3.98 1.90 3.98 3.36 5.38 3.36 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 7.68 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.54 1.20 4.54
                 1.20 4.86 6.44 4.86 6.44 4.22 6.76 4.22 6.76 4.86 7.68 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  0.88 1.22 7.46 1.54 ;
        POLYGON  7.46 4.54 7.14 4.54 7.14 3.90 6.06 3.90 6.06 4.54 4.36 4.54
                 4.36 4.22 5.74 4.22 5.74 3.58 7.46 3.58 ;
        POLYGON  3.28 4.54 1.58 4.54 1.58 4.22 0.50 4.22 0.50 4.54 0.18 4.54
                 0.18 3.58 0.50 3.58 0.50 3.90 1.58 3.90 1.58 3.58 1.90 3.58
                 1.90 4.22 3.28 4.22 ;
    END
END oai22_4

MACRO oai22_2
    CLASS CORE ;
    FOREIGN oai22_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.40 4.32 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.40 3.04 3.04 ;
        END
    END b
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.62 1.76 3.26 ;
        END
    END d
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.62 0.48 3.26 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.21  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  2.58 4.54 2.26 4.54 2.26 3.68 2.08 3.68 2.08 2.22 1.20 2.22
                 1.20 1.90 2.40 1.90 2.40 3.36 2.58 3.36 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 5.12 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.54 1.20 4.54
                 1.20 4.86 3.64 4.86 3.64 4.22 3.96 4.22 3.96 4.86 5.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  0.42 1.22 4.66 1.54 ;
        POLYGON  4.66 4.54 4.34 4.54 4.34 3.90 3.28 3.90 3.28 4.54 2.96 4.54
                 2.96 3.58 4.66 3.58 ;
        POLYGON  1.88 4.54 1.56 4.54 1.56 4.22 0.18 4.22 0.18 3.90 1.70 3.90
                 1.88 4.08 ;
    END
END oai22_2

MACRO oai22_1
    CLASS CORE ;
    FOREIGN oai22_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.68 2.72 4.32 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.36 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.80 3.04 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.72 1.76 3.04 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.69  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  2.58 4.54 2.26 4.54 2.26 3.68 2.08 3.68 2.08 2.22 1.20 2.22
                 1.20 1.90 2.40 1.90 2.40 3.36 2.58 3.36 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 5.12 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.54 1.20 4.54
                 1.20 4.86 5.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  0.42 1.22 4.66 1.54 ;
        RECT  2.96 4.22 4.66 4.54 ;
        POLYGON  1.88 4.54 1.56 4.54 1.56 4.22 0.18 4.22 0.18 3.90 1.70 3.90
                 1.88 4.08 ;
    END
END oai22_1

MACRO oai222_4
    CLASS CORE ;
    FOREIGN oai222_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.52 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.62 4.96 3.26 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.62 6.88 3.26 ;
        END
    END d
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  9.76 2.62 10.08 3.26 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  7.84 2.62 8.16 3.26 ;
        END
    END b
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.62 3.04 3.26 ;
        END
    END e
    PIN f
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.62 1.12 3.26 ;
        END
    END f
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 7.26  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.86 3.90 7.46 3.90 7.46 4.54 7.14 4.54 7.14 3.90 0.50 3.90
                 0.50 4.54 0.18 4.54 0.18 3.58 1.44 3.58 1.44 2.22 0.18 2.22
                 0.18 1.22 0.50 1.22 0.50 1.90 3.30 1.90 3.30 2.22 1.76 2.22
                 1.76 3.58 8.86 3.58 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 11.52 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  11.52 6.66 0.00 6.66 0.00 4.86 3.66 4.86 3.66 4.22 3.98 4.22
                 3.98 4.86 9.92 4.86 9.92 4.22 10.24 4.22 10.24 4.86 11.52 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  10.94 1.54 8.14 1.54 8.14 2.22 3.66 2.22 3.66 1.90 7.82 1.90
                 7.82 1.22 10.94 1.22 ;
        POLYGON  10.94 4.54 10.62 4.54 10.62 3.90 9.54 3.90 9.54 4.54 7.84 4.54
                 7.84 4.22 9.22 4.22 9.22 3.58 10.94 3.58 ;
        RECT  0.88 1.22 7.46 1.54 ;
        RECT  4.36 4.22 6.76 4.54 ;
        RECT  0.88 4.22 3.28 4.54 ;
    END
END oai222_4

MACRO oai222_2
    CLASS CORE ;
    FOREIGN oai222_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.04 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.92 2.62 6.24 3.26 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.62 4.96 3.26 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.62 3.04 3.26 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.62 4.32 3.26 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.62 2.40 3.26 ;
        END
    END e
    PIN f
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.62 0.48 3.26 ;
        END
    END f
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.66 4.54 4.34 4.54 4.34 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 3.58 0.80 3.58 0.80 1.90 1.52 1.90 1.52 2.22 1.12 2.22
                 1.12 3.58 4.66 3.58 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 7.04 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.04 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.22 2.58 4.22
                 2.58 4.86 5.72 4.86 5.72 4.22 6.04 4.22 6.04 4.86 7.04 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  6.74 4.54 6.42 4.54 6.42 3.90 5.36 3.90 5.36 4.54 5.04 4.54
                 5.04 3.58 6.74 3.58 ;
        POLYGON  6.62 1.54 5.22 1.54 5.22 2.22 3.44 2.22 3.44 1.90 4.90 1.90
                 4.90 1.22 6.62 1.22 ;
        RECT  0.42 1.22 4.54 1.54 ;
        RECT  2.96 4.22 3.96 4.54 ;
        RECT  0.88 4.22 1.88 4.54 ;
    END
END oai222_2

MACRO oai222_1
    CLASS CORE ;
    FOREIGN oai222_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.04 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.92 2.72 6.56 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.72 5.28 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.36 3.04 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.68 2.72 4.32 3.04 ;
        END
    END d
    PIN f
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.80 3.04 ;
        END
    END f
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.72 1.76 3.04 ;
        END
    END e
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.39  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.66 4.54 4.34 4.54 4.34 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 3.58 2.08 3.58 2.08 2.22 1.20 2.22 1.20 1.90 2.40 1.90
                 2.40 3.58 4.66 3.58 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 7.04 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.04 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.22 2.58 4.22
                 2.58 4.86 7.04 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  5.04 4.22 6.74 4.54 ;
        POLYGON  6.62 1.54 5.22 1.54 5.22 2.22 3.44 2.22 3.44 1.90 4.90 1.90
                 4.90 1.22 6.62 1.22 ;
        RECT  0.42 1.22 4.54 1.54 ;
        RECT  2.96 4.22 3.96 4.54 ;
        RECT  0.88 4.22 1.88 4.54 ;
    END
END oai222_1

MACRO oai221_4
    CLASS CORE ;
    FOREIGN oai221_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.24 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  8.48 2.62 8.80 3.26 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.62 6.88 3.26 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.62 3.04 3.26 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.62 0.48 3.26 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 2.62 5.60 3.26 ;
        END
    END e
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 7.26  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.46 3.90 6.06 3.90 6.06 4.54 5.74 4.54 5.74 3.90 4.66 3.90
                 4.66 4.54 4.34 4.54 4.34 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 3.58 1.62 3.58 1.62 3.04 1.44 3.04 1.44 2.72 1.62 2.72
                 1.62 2.22 0.18 2.22 0.18 1.22 0.50 1.22 0.50 1.90 3.30 1.90
                 3.30 2.22 1.94 2.22 1.94 3.58 7.46 3.58 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 10.24 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  10.24 6.66 0.00 6.66 0.00 4.86 3.66 4.86 3.66 4.22 3.98 4.22
                 3.98 4.86 5.04 4.86 5.04 4.22 5.36 4.22 5.36 4.86 8.52 4.86
                 8.52 4.22 8.84 4.22 8.84 4.86 10.24 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  4.36 1.22 9.54 1.54 ;
        POLYGON  9.54 4.54 9.22 4.54 9.22 3.90 8.14 3.90 8.14 4.54 6.44 4.54
                 6.44 4.22 7.82 4.22 7.82 3.58 9.54 3.58 ;
        POLYGON  5.38 2.22 3.66 2.22 3.66 1.54 0.88 1.54 0.88 1.22 3.98 1.22
                 3.98 1.90 5.38 1.90 ;
        RECT  0.88 4.22 3.28 4.54 ;
    END
END oai221_4

MACRO oai221_2
    CLASS CORE ;
    FOREIGN oai221_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.76 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.62 4.96 3.26 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.62 3.68 3.26 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.62 1.76 3.26 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.62 0.48 3.26 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.62 3.04 3.26 ;
        END
    END e
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.51  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.28 4.54 2.96 4.54 2.96 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 3.58 2.08 3.58 2.08 2.22 0.18 2.22 0.18 1.22 0.50 1.22
                 0.50 1.90 2.40 1.90 2.40 3.58 3.28 3.58 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 5.76 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.76 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.22 2.58 4.22
                 2.58 4.86 4.34 4.86 4.34 4.22 4.66 4.22 4.66 4.86 5.76 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  2.96 1.22 5.36 1.54 ;
        POLYGON  5.36 4.54 5.04 4.54 5.04 3.90 3.98 3.90 3.98 4.54 3.66 4.54
                 3.66 3.58 5.36 3.58 ;
        RECT  0.88 1.22 2.58 1.54 ;
        RECT  0.88 4.22 1.88 4.54 ;
    END
END oai221_2

MACRO oai221_1
    CLASS CORE ;
    FOREIGN oai221_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.76 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.62 4.96 3.26 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.62 3.68 3.26 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.53  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.62 1.76 3.26 ;
        END
    END c
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.62 3.04 3.26 ;
        END
    END e
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.53  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.62 0.48 3.26 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.72  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.28 4.54 2.96 4.54 2.96 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 3.58 2.08 3.58 2.08 2.22 0.18 2.22 0.18 1.22 0.50 1.22
                 0.50 1.90 2.40 1.90 2.40 3.58 3.28 3.58 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 5.76 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.76 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.22 2.58 4.22
                 2.58 4.86 5.76 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  2.96 1.22 5.36 1.54 ;
        RECT  3.66 4.22 5.36 4.54 ;
        RECT  0.88 1.22 2.58 1.54 ;
        RECT  0.88 4.22 1.88 4.54 ;
    END
END oai221_1

MACRO oai21_4
    CLASS CORE ;
    FOREIGN oai21_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.54 3.04 3.18 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.54 0.48 3.18 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.54 4.96 3.18 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  6.24 3.68 6.06 3.68 6.06 4.54 5.74 4.54 5.74 3.90 4.66 3.90
                 4.66 4.54 4.34 4.54 4.34 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 3.58 2.08 3.58 2.08 2.22 0.18 2.22 0.18 1.22 0.50 1.22
                 0.50 1.90 3.98 1.90 3.98 2.22 2.40 2.22 2.40 3.58 5.74 3.58
                 5.74 3.36 6.24 3.36 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 0.90 5.36 0.90 5.36 1.54 5.04 1.54 5.04 0.90 0.00 0.90
                 0.00 -0.90 6.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 6.66 0.00 6.66 0.00 4.86 5.04 4.86 5.04 4.22 5.36 4.22
                 5.36 4.86 6.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  6.06 2.22 4.34 2.22 4.34 1.54 0.88 1.54 0.88 1.22 4.66 1.22
                 4.66 1.90 5.74 1.90 5.74 1.22 6.06 1.22 ;
        RECT  0.88 4.22 3.98 4.54 ;
    END
END oai21_4

MACRO oai21_2
    CLASS CORE ;
    FOREIGN oai21_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.84 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.54 1.76 3.18 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.54 0.48 3.18 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.40 3.04 3.04 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.68 3.68 3.28 3.68 3.28 4.54 2.96 4.54 2.96 3.90 0.50 3.90
                 0.50 4.06 0.18 4.06 0.18 3.58 2.08 3.58 2.08 2.22 0.18 2.22
                 0.18 1.22 0.50 1.22 0.50 1.90 2.40 1.90 2.40 3.58 2.96 3.58
                 2.96 3.36 3.68 3.36 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  3.84 0.90 3.28 0.90 3.28 1.92 2.96 1.92 2.96 0.90 0.00 0.90
                 0.00 -0.90 3.84 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  3.84 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.22 2.58 4.22
                 2.58 4.86 3.84 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  0.88 1.22 2.58 1.54 ;
        RECT  0.88 4.22 1.88 4.54 ;
    END
END oai21_2

MACRO oai21_1
    CLASS CORE ;
    FOREIGN oai21_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.84 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.72 1.76 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.80 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.36 3.04 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.76  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.68 3.68 3.28 3.68 3.28 4.06 2.96 4.06 2.96 3.90 0.50 3.90
                 0.50 4.06 0.18 4.06 0.18 3.58 2.08 3.58 2.08 2.22 0.18 2.22
                 0.18 1.22 0.50 1.22 0.50 1.90 2.40 1.90 2.40 3.58 2.96 3.58
                 2.96 3.36 3.68 3.36 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  3.84 0.90 3.28 0.90 3.28 1.54 2.96 1.54 2.96 0.90 0.00 0.90
                 0.00 -0.90 3.84 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  3.84 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.22 2.58 4.22
                 2.58 4.86 3.84 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  0.88 1.22 2.58 1.54 ;
        RECT  0.88 4.22 1.88 4.54 ;
    END
END oai21_1

MACRO oai211_4
    CLASS CORE ;
    FOREIGN oai211_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.62 3.04 3.26 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.62 1.12 3.26 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.62 4.96 3.26 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.62 6.88 3.26 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 7.26  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.46 4.54 7.14 4.54 7.14 3.90 6.06 3.90 6.06 4.54 5.74 4.54
                 5.74 3.90 4.68 3.90 4.68 4.54 4.36 4.54 4.36 3.90 0.50 3.90
                 0.50 4.54 0.18 4.54 0.18 3.58 1.44 3.58 1.44 2.22 0.18 2.22
                 0.18 1.22 0.50 1.22 0.50 1.90 3.30 1.90 3.30 2.22 1.76 2.22
                 1.76 3.58 7.46 3.58 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 0.90 6.76 0.90 6.76 1.54 6.44 1.54 6.44 0.90 0.00 0.90
                 0.00 -0.90 7.68 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 6.66 0.00 6.66 0.00 4.86 3.66 4.86 3.66 4.22 3.98 4.22
                 3.98 4.86 5.06 4.86 5.06 4.22 5.38 4.22 5.38 4.86 6.44 4.86
                 6.44 4.22 6.76 4.22 6.76 4.86 7.68 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  7.46 2.22 5.74 2.22 5.74 1.54 4.36 1.54 4.36 1.22 6.06 1.22
                 6.06 1.90 7.46 1.90 ;
        POLYGON  5.38 2.22 3.66 2.22 3.66 1.54 0.88 1.54 0.88 1.22 3.98 1.22
                 3.98 1.90 5.38 1.90 ;
        RECT  0.88 4.22 3.28 4.54 ;
    END
END oai211_4

MACRO oai211_2
    CLASS CORE ;
    FOREIGN oai211_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.62 1.76 3.26 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.62 0.48 3.26 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.62 3.04 3.26 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.62 4.32 3.26 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.31  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.66 4.54 4.34 4.54 4.34 3.90 3.28 3.90 3.28 4.54 2.96 4.54
                 2.96 3.90 0.50 3.90 0.50 4.54 0.18 4.54 0.18 3.58 2.08 3.58
                 2.08 2.22 0.18 2.22 0.18 1.22 0.50 1.22 0.50 1.90 2.40 1.90
                 2.40 3.58 4.66 3.58 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 5.12 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.22 2.58 4.22
                 2.58 4.86 3.64 4.86 3.64 4.22 3.96 4.22 3.96 4.86 5.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  2.96 1.22 4.66 1.54 ;
        RECT  0.88 1.22 2.58 1.54 ;
        RECT  0.88 4.22 1.88 4.54 ;
    END
END oai211_2

MACRO oai211_1
    CLASS CORE ;
    FOREIGN oai211_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.72 1.76 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.80 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.36 3.04 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.72 4.64 3.04 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.47  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.66 4.54 2.96 4.54 2.96 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 3.58 2.08 3.58 2.08 2.22 0.18 2.22 0.18 1.22 0.50 1.22
                 0.50 1.90 2.40 1.90 2.40 3.58 3.28 3.58 3.28 4.22 4.66 4.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 5.12 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.22 2.58 4.22
                 2.58 4.86 5.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  2.96 1.22 4.66 1.54 ;
        RECT  0.88 1.22 2.58 1.54 ;
        RECT  0.88 4.22 1.88 4.54 ;
    END
END oai211_1

MACRO oa33_4
    CLASS CORE ;
    FOREIGN oa33_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.96 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.72 6.88 3.36 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 2.72 5.60 3.36 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.72 4.64 3.04 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.72 1.12 3.36 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.72 2.40 3.36 ;
        END
    END e
    PIN f
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.04 3.36 ;
        END
    END f
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.80 3.04 8.76 3.04 8.76 3.90 8.36 3.90 8.36 4.54 8.04 4.54
                 8.04 3.58 8.44 3.58 8.44 1.54 8.04 1.54 8.04 1.22 8.76 1.22
                 8.76 2.72 8.80 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.96 0.90 7.50 0.90 7.50 1.54 7.18 1.54 7.18 0.90 0.00 0.90
                 0.00 -0.90 8.96 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  8.96 6.66 0.00 6.66 0.00 4.86 7.23 4.86 7.23 4.22 7.55 4.22
                 7.55 4.86 8.96 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  7.96 2.44 7.64 2.44 7.64 2.40 3.68 2.40 3.68 3.52 3.96 3.52
                 3.96 4.54 3.64 4.54 3.64 3.84 3.36 3.84 3.36 2.40 0.46 2.40
                 0.46 1.22 0.78 1.22 0.78 2.08 2.62 2.08 2.62 1.86 2.94 1.86
                 2.94 2.08 7.96 2.08 ;
        RECT  1.16 1.22 6.72 1.54 ;
        RECT  5.72 4.22 6.72 4.54 ;
        RECT  4.34 4.22 5.34 4.54 ;
        RECT  2.26 4.22 3.26 4.54 ;
        RECT  0.18 4.22 1.88 4.54 ;
    END
END oa33_4

MACRO oa33_2
    CLASS CORE ;
    FOREIGN oa33_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.96 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.72 6.88 3.36 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 2.72 5.60 3.36 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.72 4.64 3.04 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.72 1.12 3.36 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.72 2.40 3.36 ;
        END
    END e
    PIN f
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.04 3.36 ;
        END
    END f
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.80 3.04 8.76 3.04 8.76 4.54 8.04 4.54 8.04 4.22 8.44 4.22
                 8.44 1.54 8.04 1.54 8.04 1.22 8.76 1.22 8.76 2.72 8.80 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.96 0.90 7.54 0.90 7.54 1.66 7.22 1.66 7.22 0.90 0.00 0.90
                 0.00 -0.90 8.96 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  8.96 6.66 0.00 6.66 0.00 4.86 7.23 4.86 7.23 4.22 7.55 4.22
                 7.55 4.86 8.96 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  7.96 2.44 7.64 2.44 7.64 2.40 3.68 2.40 3.68 3.52 3.96 3.52
                 3.96 4.54 3.64 4.54 3.64 3.84 3.36 3.84 3.36 2.40 0.46 2.40
                 0.46 1.22 0.78 1.22 0.78 2.08 2.62 2.08 2.62 1.86 2.94 1.86
                 2.94 2.08 7.96 2.08 ;
        RECT  1.16 1.22 6.72 1.54 ;
        RECT  5.72 4.22 6.72 4.54 ;
        RECT  4.34 4.22 5.34 4.54 ;
        RECT  2.26 4.22 3.26 4.54 ;
        RECT  0.18 4.22 1.88 4.54 ;
    END
END oa33_2

MACRO oa33_1
    CLASS CORE ;
    FOREIGN oa33_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.96 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.72 6.88 3.36 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 2.72 5.60 3.36 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.72 4.64 3.04 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.72 1.12 3.36 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.72 2.40 3.36 ;
        END
    END e
    PIN f
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.04 3.36 ;
        END
    END f
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.80 3.04 8.76 3.04 8.76 4.54 8.04 4.54 8.04 4.22 8.44 4.22
                 8.44 1.54 8.04 1.54 8.04 1.22 8.76 1.22 8.76 2.72 8.80 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.96 0.90 7.54 0.90 7.54 1.66 7.22 1.66 7.22 0.90 0.00 0.90
                 0.00 -0.90 8.96 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  8.96 6.66 0.00 6.66 0.00 4.86 7.26 4.86 7.26 3.98 7.58 3.98
                 7.58 4.86 8.96 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  7.96 2.44 7.64 2.44 7.64 2.40 3.68 2.40 3.68 3.52 3.96 3.52
                 3.96 4.54 3.64 4.54 3.64 3.84 3.36 3.84 3.36 2.40 0.46 2.40
                 0.46 1.22 0.78 1.22 0.78 2.08 2.62 2.08 2.62 1.86 2.94 1.86
                 2.94 2.08 7.96 2.08 ;
        RECT  1.16 1.22 6.72 1.54 ;
        RECT  5.72 4.22 6.72 4.54 ;
        RECT  4.34 4.22 5.34 4.54 ;
        RECT  2.26 4.22 3.26 4.54 ;
        RECT  0.18 4.22 1.88 4.54 ;
    END
END oa33_1

MACRO oa32_4
    CLASS CORE ;
    FOREIGN oa32_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 2.72 5.60 3.36 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.94 2.72 4.32 3.36 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.04 3.36 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.72 1.12 3.36 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.72 1.76 3.36 ;
        END
    END e
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.52 3.04 7.38 3.04 7.38 3.42 6.98 3.42 6.98 4.54 6.66 4.54
                 6.66 3.10 7.06 3.10 7.06 1.54 6.66 1.54 6.66 1.22 7.38 1.22
                 7.38 2.72 7.52 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 0.90 6.12 0.90 6.12 1.54 5.80 1.54 5.80 0.90 0.00 0.90
                 0.00 -0.90 7.68 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 6.66 0.00 6.66 0.00 4.86 5.85 4.86 5.85 4.22 6.17 4.22
                 6.17 4.86 7.68 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  6.58 2.44 6.26 2.44 6.26 2.40 2.40 2.40 2.40 3.65 2.58 3.65
                 2.58 4.54 2.26 4.54 2.26 3.94 2.08 3.94 2.08 2.40 1.24 2.40
                 1.24 1.86 1.56 1.86 1.56 2.08 6.58 2.08 ;
        RECT  0.46 1.22 5.34 1.54 ;
        RECT  4.34 4.22 5.34 4.54 ;
        RECT  2.96 4.22 3.96 4.54 ;
        RECT  0.18 4.22 1.88 4.54 ;
    END
END oa32_4

MACRO oa32_2
    CLASS CORE ;
    FOREIGN oa32_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 2.72 5.60 3.36 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.94 2.72 4.32 3.36 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.04 3.36 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.72 1.12 3.36 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.72 1.76 3.36 ;
        END
    END e
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.52 3.04 7.38 3.04 7.38 4.54 6.66 4.54 6.66 4.22 7.06 4.22
                 7.06 1.54 6.66 1.54 6.66 1.22 7.38 1.22 7.38 2.72 7.52 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 0.90 6.16 0.90 6.16 1.66 5.84 1.66 5.84 0.90 0.00 0.90
                 0.00 -0.90 7.68 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 6.66 0.00 6.66 0.00 4.86 5.85 4.86 5.85 4.22 6.17 4.22
                 6.17 4.86 7.68 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  6.58 2.44 6.26 2.44 6.26 2.40 2.40 2.40 2.40 3.65 2.58 3.65
                 2.58 4.54 2.26 4.54 2.26 3.94 2.08 3.94 2.08 2.40 1.24 2.40
                 1.24 1.86 1.56 1.86 1.56 2.08 6.58 2.08 ;
        RECT  0.46 1.22 5.34 1.54 ;
        RECT  4.34 4.22 5.34 4.54 ;
        RECT  2.96 4.22 3.96 4.54 ;
        RECT  0.18 4.22 1.88 4.54 ;
    END
END oa32_2

MACRO oa32_1
    CLASS CORE ;
    FOREIGN oa32_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 2.72 5.60 3.36 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.94 2.72 4.32 3.36 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.04 3.36 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.72 1.12 3.36 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.72 1.76 3.36 ;
        END
    END e
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.52 3.04 7.38 3.04 7.38 4.54 6.66 4.54 6.66 4.22 7.06 4.22
                 7.06 1.54 6.66 1.54 6.66 1.22 7.38 1.22 7.38 2.72 7.52 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 0.90 6.16 0.90 6.16 1.66 5.84 1.66 5.84 0.90 0.00 0.90
                 0.00 -0.90 7.68 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 6.66 0.00 6.66 0.00 4.86 5.88 4.86 5.88 3.98 6.20 3.98
                 6.20 4.86 7.68 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  6.58 2.44 6.26 2.44 6.26 2.40 2.40 2.40 2.40 3.65 2.58 3.65
                 2.58 4.54 2.26 4.54 2.26 3.94 2.08 3.94 2.08 2.40 1.24 2.40
                 1.24 1.86 1.56 1.86 1.56 2.08 6.58 2.08 ;
        RECT  0.46 1.22 5.34 1.54 ;
        RECT  4.34 4.22 5.34 4.54 ;
        RECT  2.96 4.22 3.96 4.54 ;
        RECT  0.18 4.22 1.88 4.54 ;
    END
END oa32_1

MACRO oa31_4
    CLASS CORE ;
    FOREIGN oa31_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.72 4.32 3.36 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.04 3.36 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.72 1.76 3.36 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.72 1.12 3.36 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  6.24 3.42 5.84 3.42 5.84 4.54 5.52 4.54 5.52 3.10 5.92 3.10
                 5.92 1.54 5.52 1.54 5.52 1.22 6.24 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 0.90 5.02 0.90 5.02 1.54 4.70 1.54 4.70 0.90 0.00 0.90
                 0.00 -0.90 6.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 6.66 0.00 6.66 0.00 4.86 0.42 4.86 0.42 4.38 0.74 4.38
                 0.74 4.86 4.71 4.86 4.71 4.22 5.03 4.22 5.03 4.86 6.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  5.44 2.44 5.12 2.44 5.12 2.40 0.48 2.40 0.48 3.74 1.44 3.74
                 1.44 4.06 0.16 4.06 0.16 1.34 0.50 1.34 0.50 1.66 0.48 1.66
                 0.48 2.08 5.44 2.08 ;
        RECT  0.88 1.22 4.20 1.54 ;
        RECT  3.20 4.22 4.20 4.54 ;
        RECT  1.82 4.22 2.82 4.54 ;
    END
END oa31_4

MACRO oa31_2
    CLASS CORE ;
    FOREIGN oa31_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.72 4.32 3.36 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.04 3.36 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.72 1.76 3.36 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.72 1.12 3.36 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  6.24 4.54 5.52 4.54 5.52 4.22 5.92 4.22 5.92 1.54 5.52 1.54
                 5.52 1.22 6.24 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 0.90 5.02 0.90 5.02 1.20 4.70 1.20 4.70 0.90 0.00 0.90
                 0.00 -0.90 6.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 6.66 0.00 6.66 0.00 4.86 0.42 4.86 0.42 4.38 0.74 4.38
                 0.74 4.86 4.71 4.86 4.71 4.22 5.03 4.22 5.03 4.86 6.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  5.44 2.44 5.12 2.44 5.12 2.40 0.48 2.40 0.48 3.74 1.44 3.74
                 1.44 4.06 0.16 4.06 0.16 1.34 0.50 1.34 0.50 1.66 0.48 1.66
                 0.48 2.08 5.44 2.08 ;
        RECT  0.88 1.22 4.20 1.54 ;
        RECT  3.20 4.22 4.20 4.54 ;
        RECT  1.82 4.22 2.82 4.54 ;
    END
END oa31_2

MACRO oa31_1
    CLASS CORE ;
    FOREIGN oa31_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.72 4.32 3.36 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.04 3.36 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.72 1.76 3.36 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.72 1.12 3.36 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  6.24 4.54 5.52 4.54 5.52 4.22 5.92 4.22 5.92 1.54 5.52 1.54
                 5.52 1.22 6.24 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 0.90 5.02 0.90 5.02 1.66 4.70 1.66 4.70 0.90 0.00 0.90
                 0.00 -0.90 6.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 6.66 0.00 6.66 0.00 4.86 4.74 4.86 4.74 3.98 5.06 3.98
                 5.06 4.86 6.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  5.44 2.44 5.12 2.44 5.12 2.40 0.48 2.40 0.48 3.74 1.44 3.74
                 1.44 4.06 0.16 4.06 0.16 1.34 0.50 1.34 0.50 1.66 0.48 1.66
                 0.48 2.08 5.44 2.08 ;
        RECT  0.88 1.22 4.20 1.54 ;
        RECT  3.20 4.22 4.20 4.54 ;
        RECT  1.82 4.22 2.82 4.54 ;
    END
END oa31_1

MACRO oa22_4
    CLASS CORE ;
    FOREIGN oa22_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.68 2.72 4.32 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.36 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.80 3.04 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.72 1.76 3.04 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  6.24 3.04 6.04 3.04 6.04 4.54 5.72 4.54 5.72 1.64 6.04 1.64
                 6.04 2.72 6.24 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 0.90 5.34 0.90 5.34 1.54 5.02 1.54 5.02 0.90 0.00 0.90
                 0.00 -0.90 6.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.54 1.20 4.54
                 1.20 4.86 5.02 4.86 5.02 3.66 5.34 3.66 5.34 4.86 6.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  5.40 2.44 5.08 2.44 5.08 2.40 2.40 2.40 2.40 3.33 2.58 3.33
                 2.58 4.54 2.26 4.54 2.26 3.65 2.08 3.65 2.08 2.22 1.20 2.22
                 1.20 1.90 2.40 1.90 2.40 2.08 5.40 2.08 ;
        RECT  0.42 1.22 4.66 1.54 ;
        RECT  2.96 4.22 4.66 4.54 ;
        POLYGON  1.88 4.54 1.56 4.54 1.56 4.22 0.18 4.22 0.18 3.90 1.88 3.90 ;
    END
END oa22_4

MACRO oa22_2
    CLASS CORE ;
    FOREIGN oa22_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.68 2.72 4.32 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.36 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.80 3.04 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.72 1.76 3.04 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  6.24 3.04 6.04 3.04 6.04 4.06 5.72 4.06 5.72 1.64 6.04 1.64
                 6.04 2.72 6.24 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 0.90 5.34 0.90 5.34 1.54 5.02 1.54 5.02 0.90 0.00 0.90
                 0.00 -0.90 6.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.54 1.20 4.54
                 1.20 4.86 5.02 4.86 5.02 4.22 5.34 4.22 5.34 4.86 6.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  5.40 2.44 5.08 2.44 5.08 2.40 2.40 2.40 2.40 3.33 2.58 3.33
                 2.58 4.54 2.26 4.54 2.26 3.65 2.08 3.65 2.08 2.22 1.20 2.22
                 1.20 1.90 2.40 1.90 2.40 2.08 5.40 2.08 ;
        RECT  0.42 1.22 4.66 1.54 ;
        RECT  2.96 4.22 4.66 4.54 ;
        POLYGON  1.88 4.54 1.56 4.54 1.56 4.22 0.18 4.22 0.18 3.90 1.88 3.90 ;
    END
END oa22_2

MACRO oa22_1
    CLASS CORE ;
    FOREIGN oa22_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.68 2.72 4.32 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.36 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.80 3.04 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.72 1.76 3.04 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  6.24 3.04 6.04 3.04 6.04 4.30 5.72 4.30 5.72 1.64 6.04 1.64
                 6.04 2.72 6.24 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 0.90 5.34 0.90 5.34 1.20 5.02 1.20 5.02 0.90 0.00 0.90
                 0.00 -0.90 6.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.54 1.20 4.54
                 1.20 4.86 5.02 4.86 5.02 4.28 5.34 4.28 5.34 4.86 6.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  5.40 2.44 5.08 2.44 5.08 2.40 2.40 2.40 2.40 3.33 2.58 3.33
                 2.58 4.54 2.26 4.54 2.26 3.65 2.08 3.65 2.08 2.22 1.20 2.22
                 1.20 1.90 2.40 1.90 2.40 2.08 5.40 2.08 ;
        RECT  0.42 1.22 4.66 1.54 ;
        RECT  2.96 4.22 4.66 4.54 ;
        POLYGON  1.88 4.54 1.56 4.54 1.56 4.22 0.18 4.22 0.18 3.90 1.88 3.90 ;
    END
END oa22_1

MACRO oa222_4
    CLASS CORE ;
    FOREIGN oa222_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.32 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.92 2.40 6.24 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.72 5.28 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.36 3.04 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.68 2.72 4.32 3.04 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.72 1.76 3.04 ;
        END
    END e
    PIN f
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.80 3.04 ;
        END
    END f
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.16 3.04 8.00 3.04 8.00 3.42 7.68 3.42 7.68 4.54 7.36 4.54
                 7.36 3.10 7.68 3.10 7.68 1.22 8.00 1.22 8.00 2.72 8.16 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 0.90 7.30 0.90 7.30 1.54 6.98 1.54 6.98 0.90 0.00 0.90
                 0.00 -0.90 8.32 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.22 2.58 4.22
                 2.58 4.86 6.54 4.86 6.54 4.22 6.86 4.22 6.86 4.86 8.32 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  7.04 3.90 4.66 3.90 4.66 4.54 4.34 4.54 4.34 3.90 0.50 3.90
                 0.50 4.54 0.18 4.54 0.18 3.58 2.08 3.58 2.08 2.22 1.20 2.22
                 1.20 1.90 2.40 1.90 2.40 3.58 6.72 3.58 6.72 2.12 7.04 2.12 ;
        POLYGON  6.62 1.54 5.22 1.54 5.22 2.22 3.44 2.22 3.44 1.90 4.90 1.90
                 4.90 1.22 6.62 1.22 ;
        RECT  5.04 4.22 6.04 4.54 ;
        RECT  0.42 1.22 4.54 1.54 ;
        RECT  2.96 4.22 3.96 4.54 ;
        RECT  0.88 4.22 1.88 4.54 ;
    END
END oa222_4

MACRO oa222_2
    CLASS CORE ;
    FOREIGN oa222_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.32 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.92 2.72 6.56 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.72 5.28 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.36 3.04 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.68 2.72 4.32 3.04 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.72 1.76 3.04 ;
        END
    END e
    PIN f
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.80 3.04 ;
        END
    END f
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.16 3.04 8.00 3.04 8.00 4.54 7.36 4.54 7.36 4.22 7.68 4.22
                 7.68 1.22 8.00 1.22 8.00 2.72 8.16 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 0.90 7.30 0.90 7.30 1.54 6.98 1.54 6.98 0.90 0.00 0.90
                 0.00 -0.90 8.32 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.22 2.58 4.22
                 2.58 4.86 6.54 4.86 6.54 4.22 6.86 4.22 6.86 4.86 8.32 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  7.35 3.90 4.66 3.90 4.66 4.54 4.34 4.54 4.34 3.90 0.50 3.90
                 0.50 4.54 0.18 4.54 0.18 3.58 2.08 3.58 2.08 2.22 1.20 2.22
                 1.20 1.90 2.40 1.90 2.40 3.58 7.03 3.58 7.03 2.12 7.35 2.12 ;
        POLYGON  6.62 1.54 5.22 1.54 5.22 2.22 3.44 2.22 3.44 1.90 4.90 1.90
                 4.90 1.22 6.62 1.22 ;
        RECT  5.04 4.22 6.04 4.54 ;
        RECT  0.42 1.22 4.54 1.54 ;
        RECT  2.96 4.22 3.96 4.54 ;
        RECT  0.88 4.22 1.88 4.54 ;
    END
END oa222_2

MACRO oa222_1
    CLASS CORE ;
    FOREIGN oa222_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.32 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.92 2.72 6.56 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.72 5.28 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.36 3.04 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.68 2.72 4.32 3.04 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.72 1.76 3.04 ;
        END
    END e
    PIN f
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.80 3.04 ;
        END
    END f
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.16 3.04 8.00 3.04 8.00 4.54 7.36 4.54 7.36 4.22 7.68 4.22
                 7.68 1.22 8.00 1.22 8.00 2.72 8.16 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 0.90 7.30 0.90 7.30 1.54 6.98 1.54 6.98 0.90 0.00 0.90
                 0.00 -0.90 8.32 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.22 2.58 4.22
                 2.58 4.86 6.53 4.86 6.53 4.28 6.85 4.28 6.85 4.86 8.32 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  7.35 3.90 4.66 3.90 4.66 4.54 4.34 4.54 4.34 3.90 0.50 3.90
                 0.50 4.54 0.18 4.54 0.18 3.58 2.08 3.58 2.08 2.22 1.20 2.22
                 1.20 1.90 2.40 1.90 2.40 3.58 7.03 3.58 7.03 2.12 7.35 2.12 ;
        POLYGON  6.62 1.54 5.22 1.54 5.22 2.22 3.44 2.22 3.44 1.90 4.90 1.90
                 4.90 1.22 6.62 1.22 ;
        RECT  5.04 4.22 6.04 4.54 ;
        RECT  0.42 1.22 4.54 1.54 ;
        RECT  2.96 4.22 3.96 4.54 ;
        RECT  0.88 4.22 1.88 4.54 ;
    END
END oa222_1

MACRO oa221_4
    CLASS CORE ;
    FOREIGN oa221_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.96 2.72 5.60 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.68 2.72 4.32 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.72 1.76 3.04 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.80 3.04 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.36 3.04 ;
        END
    END e
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.52 3.04 7.14 3.04 7.14 4.54 6.82 4.54 6.82 1.22 7.14 1.22
                 7.14 2.72 7.52 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 0.90 6.44 0.90 6.44 1.54 6.12 1.54 6.12 0.90 0.00 0.90
                 0.00 -0.90 7.68 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 6.66 0.00 6.66 0.00 4.86 2.46 4.86 2.46 4.22 2.78 4.22
                 2.78 4.86 5.44 4.86 5.44 4.22 5.76 4.22 5.76 4.86 6.12 4.86
                 6.12 3.66 6.44 3.66 6.44 4.86 7.68 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  6.49 2.44 6.17 2.44 6.17 2.40 2.40 2.40 2.40 3.58 3.68 3.58
                 3.68 4.54 3.36 4.54 3.36 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 3.58 2.08 3.58 2.08 2.22 1.20 2.22 1.20 1.90 2.40 1.90
                 2.40 2.08 6.49 2.08 ;
        RECT  3.36 1.22 5.76 1.54 ;
        RECT  4.06 4.22 5.06 4.54 ;
        RECT  0.42 1.22 2.98 1.54 ;
        RECT  0.88 4.22 1.88 4.54 ;
    END
END oa221_4

MACRO oa221_2
    CLASS CORE ;
    FOREIGN oa221_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.96 2.72 5.60 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.68 2.72 4.32 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.72 1.76 3.04 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.80 3.04 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.36 3.04 ;
        END
    END e
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.52 3.04 7.14 3.04 7.14 4.54 6.82 4.54 6.82 1.22 7.14 1.22
                 7.14 2.72 7.52 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 0.90 6.44 0.90 6.44 1.54 6.12 1.54 6.12 0.90 0.00 0.90
                 0.00 -0.90 7.68 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 6.66 0.00 6.66 0.00 4.86 2.46 4.86 2.46 4.22 2.78 4.22
                 2.78 4.86 5.44 4.86 5.44 4.22 6.44 4.22 6.44 4.86 7.68 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  6.49 2.44 6.17 2.44 6.17 2.40 2.40 2.40 2.40 3.58 3.68 3.58
                 3.68 4.54 3.36 4.54 3.36 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 3.58 2.08 3.58 2.08 2.22 1.20 2.22 1.20 1.90 2.40 1.90
                 2.40 2.08 6.49 2.08 ;
        RECT  3.36 1.22 5.76 1.54 ;
        RECT  4.06 4.22 5.06 4.54 ;
        RECT  0.42 1.22 2.98 1.54 ;
        RECT  0.88 4.22 1.88 4.54 ;
    END
END oa221_2

MACRO oa221_1
    CLASS CORE ;
    FOREIGN oa221_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.04 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.96 2.72 5.60 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.72 4.64 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 3.26 2.08 3.68 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 3.26 1.12 3.90 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.72 3.04 3.04 ;
        END
    END e
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  6.88 3.04 6.74 3.04 6.74 4.54 6.42 4.54 6.42 1.22 6.74 1.22
                 6.74 2.72 6.88 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  7.04 0.90 6.04 0.90 6.04 1.66 5.72 1.66 5.72 0.90 0.00 0.90
                 0.00 -0.90 7.04 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.04 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.22 2.58 4.22
                 2.58 4.86 5.04 4.86 5.04 4.22 5.36 4.22 5.36 4.86 5.72 4.86
                 5.72 4.28 6.04 4.28 6.04 4.86 7.04 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  6.10 2.44 5.78 2.44 5.78 2.40 3.68 2.40 3.68 3.68 3.28 3.68
                 3.28 4.54 2.96 4.54 2.96 3.36 3.36 3.36 3.36 2.40 0.48 2.40
                 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54 0.16 1.90 0.50 1.90
                 0.50 2.08 1.58 2.08 1.58 1.90 1.90 1.90 1.90 2.08 6.10 2.08 ;
        RECT  2.96 1.22 5.36 1.54 ;
        RECT  3.66 4.22 4.66 4.54 ;
        POLYGON  2.58 1.54 1.20 1.54 1.20 1.76 0.88 1.76 0.88 1.22 2.58 1.22 ;
        RECT  0.88 4.22 1.88 4.54 ;
    END
END oa221_1

MACRO oa21_4
    CLASS CORE ;
    FOREIGN oa21_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.72 1.76 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.80 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.36 3.04 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.96 3.42 4.66 3.42 4.66 4.54 4.34 4.54 4.34 3.10 4.64 3.10
                 4.64 1.54 4.34 1.54 4.34 1.22 4.96 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 0.90 3.82 0.90 3.82 1.54 3.50 1.54 3.50 0.90 0.00 0.90
                 0.00 -0.90 5.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.22 2.58 4.22
                 2.58 4.86 3.64 4.86 3.64 3.66 3.96 3.66 3.96 4.86 5.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.32 2.44 4.00 2.44 4.00 2.40 2.40 2.40 2.40 3.58 3.28 3.58
                 3.28 4.06 2.96 4.06 2.96 3.90 0.50 3.90 0.50 4.06 0.18 4.06
                 0.18 3.58 2.08 3.58 2.08 2.22 1.20 2.22 1.20 1.90 2.40 1.90
                 2.40 2.08 4.32 2.08 ;
        RECT  0.42 1.22 2.98 1.54 ;
        RECT  0.88 4.22 1.88 4.54 ;
    END
END oa21_4

MACRO oa21_2
    CLASS CORE ;
    FOREIGN oa21_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.72 1.76 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.80 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.36 3.04 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.96 4.06 4.34 4.06 4.34 3.74 4.64 3.74 4.64 1.54 4.34 1.54
                 4.34 1.22 4.96 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 0.90 3.84 0.90 3.84 1.54 3.52 1.54 3.52 0.90 0.00 0.90
                 0.00 -0.90 5.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.22 2.58 4.22
                 2.58 4.86 3.64 4.86 3.64 4.42 3.96 4.42 3.96 4.86 5.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.32 2.44 4.00 2.44 4.00 2.40 2.40 2.40 2.40 3.58 3.28 3.58
                 3.28 4.06 2.96 4.06 2.96 3.90 0.50 3.90 0.50 4.06 0.18 4.06
                 0.18 3.58 2.08 3.58 2.08 2.22 1.20 2.22 1.20 1.90 2.40 1.90
                 2.40 2.08 4.32 2.08 ;
        RECT  0.42 1.22 2.98 1.54 ;
        RECT  0.88 4.22 1.88 4.54 ;
    END
END oa21_2

MACRO oa21_1
    CLASS CORE ;
    FOREIGN oa21_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.72 1.76 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.80 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.36 3.04 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.96 4.30 4.34 4.30 4.34 3.98 4.64 3.98 4.64 1.54 4.34 1.54
                 4.34 1.22 4.96 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 0.90 3.84 0.90 3.84 1.54 3.52 1.54 3.52 0.90 0.00 0.90
                 0.00 -0.90 5.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.22 2.58 4.22
                 2.58 4.86 3.64 4.86 3.64 4.42 3.96 4.42 3.96 4.86 5.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.32 2.44 4.00 2.44 4.00 2.40 2.40 2.40 2.40 3.58 3.28 3.58
                 3.28 4.06 2.96 4.06 2.96 3.90 0.50 3.90 0.50 4.06 0.18 4.06
                 0.18 3.58 2.08 3.58 2.08 2.22 1.20 2.22 1.20 1.90 2.40 1.90
                 2.40 2.08 4.32 2.08 ;
        RECT  0.42 1.22 2.98 1.54 ;
        RECT  0.88 4.22 1.88 4.54 ;
    END
END oa21_1

MACRO oa211_4
    CLASS CORE ;
    FOREIGN oa211_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.72 1.76 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.80 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.36 3.04 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.72 4.64 3.04 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  6.24 4.54 5.68 4.54 5.68 4.22 5.92 4.22 5.92 1.54 5.68 1.54
                 5.68 1.22 6.24 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 0.90 5.18 0.90 5.18 1.54 4.86 1.54 4.86 0.90 0.00 0.90
                 0.00 -0.90 6.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.22 2.58 4.22
                 2.58 4.86 4.67 4.86 4.67 4.22 4.99 4.22 4.99 4.86 6.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  5.60 2.94 4.96 2.94 4.96 2.40 2.40 2.40 2.40 3.58 3.28 3.58
                 3.28 4.22 3.96 4.22 3.96 4.54 2.96 4.54 2.96 3.90 0.50 3.90
                 0.50 4.54 0.18 4.54 0.18 3.58 2.08 3.58 2.08 2.22 1.20 2.22
                 1.20 1.90 2.40 1.90 2.40 2.08 5.28 2.08 5.28 2.62 5.60 2.62 ;
        RECT  3.36 1.22 4.36 1.54 ;
        RECT  0.42 1.22 2.98 1.54 ;
        RECT  0.88 4.22 1.88 4.54 ;
    END
END oa211_4

MACRO oa211_2
    CLASS CORE ;
    FOREIGN oa211_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.72 1.76 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.80 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.36 3.04 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.72 4.64 3.04 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  6.24 4.54 5.68 4.54 5.68 4.22 5.92 4.22 5.92 1.54 5.68 1.54
                 5.68 1.22 6.24 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 0.90 5.18 0.90 5.18 1.54 4.86 1.54 4.86 0.90 0.00 0.90
                 0.00 -0.90 6.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.22 2.58 4.22
                 2.58 4.86 4.67 4.86 4.67 4.22 4.99 4.22 4.99 4.86 6.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  5.60 3.04 4.96 3.04 4.96 2.40 2.40 2.40 2.40 3.58 3.28 3.58
                 3.28 4.22 3.96 4.22 3.96 4.54 2.96 4.54 2.96 3.90 0.50 3.90
                 0.50 4.54 0.18 4.54 0.18 3.58 2.08 3.58 2.08 2.22 1.20 2.22
                 1.20 1.90 2.40 1.90 2.40 2.08 5.28 2.08 5.28 2.72 5.60 2.72 ;
        RECT  3.36 1.22 4.36 1.54 ;
        RECT  0.42 1.22 2.98 1.54 ;
        RECT  0.88 4.22 1.88 4.54 ;
    END
END oa211_2

MACRO oa211_1
    CLASS CORE ;
    FOREIGN oa211_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.72 1.76 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.80 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.36 3.04 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.72 4.64 3.04 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  6.24 4.54 5.68 4.54 5.68 4.22 5.92 4.22 5.92 1.54 5.68 1.54
                 5.68 1.22 6.24 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 0.90 5.18 0.90 5.18 1.54 4.86 1.54 4.86 0.90 0.00 0.90
                 0.00 -0.90 6.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.22 2.58 4.22
                 2.58 4.86 4.67 4.86 4.67 4.28 4.99 4.28 4.99 4.86 6.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  5.60 3.04 4.96 3.04 4.96 2.40 2.40 2.40 2.40 3.58 3.28 3.58
                 3.28 4.22 3.96 4.22 3.96 4.54 2.96 4.54 2.96 3.90 0.50 3.90
                 0.50 4.54 0.18 4.54 0.18 3.58 2.08 3.58 2.08 2.22 1.20 2.22
                 1.20 1.90 2.40 1.90 2.40 2.08 5.28 2.08 5.28 2.72 5.60 2.72 ;
        RECT  3.36 1.22 4.36 1.54 ;
        RECT  0.42 1.22 2.98 1.54 ;
        RECT  0.88 4.22 1.88 4.54 ;
    END
END oa211_1

MACRO nor4_8
    CLASS CORE ;
    FOREIGN nor4_8 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.16 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 1.76 0.48 2.40 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 1.76 2.72 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 1.86 4.32 2.50 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.08 2.82 2.40 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.29  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  11.96 1.74 10.56 1.74 10.56 2.72 10.72 2.72 10.72 3.04
                 10.56 3.04 10.56 3.78 11.64 3.78 11.64 3.10 11.96 3.10
                 11.96 4.10 8.84 4.10 8.84 3.16 9.16 3.16 9.16 3.78 10.24 3.78
                 10.24 1.74 8.84 1.74 8.84 1.42 11.96 1.42 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  12.16 0.90 4.32 0.90 4.32 1.54 4.00 1.54 4.00 0.90 2.92 0.90
                 2.92 1.54 2.60 1.54 2.60 0.90 2.24 0.90 2.24 1.54 1.92 1.54
                 1.92 0.90 0.00 0.90 0.00 -0.90 12.16 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  12.16 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.22 2.58 4.22
                 2.58 4.86 9.54 4.86 9.54 4.42 9.86 4.42 9.86 4.86 10.94 4.86
                 10.94 4.42 11.26 4.42 11.26 4.86 12.16 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  9.78 2.44 8.48 2.44 8.48 4.54 5.02 4.54 5.02 4.22 8.16 4.22
                 8.16 2.18 6.76 2.18 6.76 1.86 8.16 1.86 8.16 1.45 8.48 1.45
                 8.48 2.12 9.78 2.12 ;
        RECT  4.68 1.22 7.78 1.54 ;
        POLYGON  7.22 3.90 0.50 3.90 0.50 4.54 0.18 4.54 0.18 3.58 0.80 3.58
                 0.80 1.22 1.54 1.22 1.54 1.54 1.12 1.54 1.12 3.58 6.90 3.58
                 6.90 2.93 7.22 2.93 ;
        POLYGON  5.43 3.26 3.30 3.26 3.30 1.22 3.62 1.22 3.62 2.94 5.43 2.94 ;
        RECT  2.96 4.22 3.96 4.54 ;
        RECT  0.88 4.22 1.88 4.54 ;
    END
END nor4_8

MACRO nor4_4
    CLASS CORE ;
    FOREIGN nor4_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.60 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 1.76 0.48 2.40 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 1.76 2.72 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 1.86 4.32 2.50 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.08 2.82 2.40 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.97  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.12 4.54 7.80 4.54 7.80 3.68 7.20 3.68 7.20 3.36 7.80 3.36
                 7.80 1.22 8.12 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  9.60 0.90 8.82 0.90 8.82 1.55 8.50 1.55 8.50 0.90 7.29 0.90
                 7.29 1.54 6.97 1.54 6.97 0.90 4.32 0.90 4.32 1.54 4.00 1.54
                 4.00 0.90 2.92 0.90 2.92 1.54 2.60 1.54 2.60 0.90 2.24 0.90
                 2.24 1.54 1.92 1.54 1.92 0.90 0.00 0.90 0.00 -0.90 9.60 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  9.60 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.22 2.58 4.22
                 2.58 4.86 5.02 4.86 5.02 4.22 5.34 4.22 5.34 4.86 7.10 4.86
                 7.10 4.22 7.42 4.22 7.42 4.86 8.50 4.86 8.50 4.20 8.82 4.20
                 8.82 4.86 9.60 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  6.98 3.01 6.60 3.01 6.60 4.54 5.72 4.54 5.72 4.22 6.28 4.22
                 6.28 2.18 4.78 2.18 4.78 1.22 5.10 1.22 5.10 1.86 6.60 1.86
                 6.60 2.69 6.98 2.69 ;
        RECT  5.48 1.22 6.48 1.54 ;
        POLYGON  5.96 2.94 5.08 2.94 5.08 3.26 3.30 3.26 3.30 1.22 3.62 1.22
                 3.62 2.94 4.76 2.94 4.76 2.62 5.96 2.62 ;
        POLYGON  5.72 3.90 0.50 3.90 0.50 4.54 0.18 4.54 0.18 3.58 0.80 3.58
                 0.80 1.22 1.54 1.22 1.54 1.54 1.12 1.54 1.12 3.58 5.40 3.58
                 5.40 3.26 5.72 3.26 ;
        RECT  2.96 4.22 3.96 4.54 ;
        RECT  0.88 4.22 1.88 4.54 ;
    END
END nor4_4

MACRO nor4_2
    CLASS CORE ;
    FOREIGN nor4_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.32 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 1.76 0.48 2.40 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 1.76 2.72 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 1.86 4.32 2.50 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.08 2.82 2.40 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.12 4.54 7.80 4.54 7.80 3.68 7.20 3.68 7.20 3.36 7.80 3.36
                 7.80 1.22 8.12 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 0.90 7.34 0.90 7.34 1.48 7.02 1.48 7.02 0.90 4.32 0.90
                 4.32 1.54 4.00 1.54 4.00 0.90 2.92 0.90 2.92 1.54 2.60 1.54
                 2.60 0.90 2.24 0.90 2.24 1.54 1.92 1.54 1.92 0.90 0.00 0.90
                 0.00 -0.90 8.32 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.22 2.58 4.22
                 2.58 4.86 5.02 4.86 5.02 4.22 5.34 4.22 5.34 4.86 7.10 4.86
                 7.10 4.22 7.42 4.22 7.42 4.86 8.32 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  6.90 2.99 6.60 2.99 6.60 4.54 5.72 4.54 5.72 4.22 6.28 4.22
                 6.28 2.18 4.78 2.18 4.78 1.22 5.10 1.22 5.10 1.86 6.60 1.86
                 6.60 2.67 6.90 2.67 ;
        RECT  5.48 1.22 6.48 1.54 ;
        POLYGON  5.96 2.94 5.08 2.94 5.08 3.26 3.30 3.26 3.30 1.22 3.62 1.22
                 3.62 2.94 4.76 2.94 4.76 2.62 5.96 2.62 ;
        POLYGON  5.72 3.90 0.50 3.90 0.50 4.54 0.18 4.54 0.18 3.58 0.80 3.58
                 0.80 1.22 1.54 1.22 1.54 1.54 1.12 1.54 1.12 3.58 5.40 3.58
                 5.40 3.26 5.72 3.26 ;
        RECT  2.96 4.22 3.96 4.54 ;
        RECT  0.88 4.22 1.88 4.54 ;
    END
END nor4_2

MACRO nor4_1
    CLASS CORE ;
    FOREIGN nor4_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.32 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 1.76 0.48 2.40 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 1.76 2.72 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 1.79 4.32 2.43 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.08 2.82 2.40 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.12 4.54 7.80 4.54 7.80 3.68 7.20 3.68 7.20 3.36 7.80 3.36
                 7.80 1.22 8.12 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 0.90 7.34 0.90 7.34 1.54 7.02 1.54 7.02 0.90 4.32 0.90
                 4.32 1.18 4.00 1.18 4.00 0.90 2.92 0.90 2.92 1.19 2.60 1.19
                 2.60 0.90 2.24 0.90 2.24 1.18 1.92 1.18 1.92 0.90 0.00 0.90
                 0.00 -0.90 8.32 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.22 2.58 4.22
                 2.58 4.86 5.02 4.86 5.02 4.22 5.34 4.22 5.34 4.86 7.10 4.86
                 7.10 4.28 7.42 4.28 7.42 4.86 8.32 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  6.90 2.99 6.60 2.99 6.60 4.54 5.72 4.54 5.72 4.22 6.28 4.22
                 6.28 2.18 4.78 2.18 4.78 1.22 5.10 1.22 5.10 1.86 6.60 1.86
                 6.60 2.67 6.90 2.67 ;
        RECT  5.48 1.22 6.48 1.54 ;
        POLYGON  5.96 2.94 5.08 2.94 5.08 3.26 3.14 3.26 3.14 1.44 3.30 1.44
                 3.30 1.22 3.62 1.22 3.62 1.76 3.46 1.76 3.46 2.94 4.76 2.94
                 4.76 2.62 5.96 2.62 ;
        POLYGON  5.72 3.90 0.50 3.90 0.50 4.54 0.18 4.54 0.18 3.58 0.80 3.58
                 0.80 1.22 1.54 1.22 1.54 1.54 1.12 1.54 1.12 3.58 5.40 3.58
                 5.40 3.26 5.72 3.26 ;
        RECT  2.96 4.22 3.96 4.54 ;
        RECT  0.88 4.22 1.88 4.54 ;
    END
END nor4_1

MACRO nor3_8
    CLASS CORE ;
    FOREIGN nor3_8 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.20 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 5.30  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  16.76 2.08 17.76 2.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 5.30  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.40 2.08 11.48 2.43 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 5.30  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.08 1.76 2.43 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 13.75  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  18.66 3.90 12.74 3.90 12.74 2.40 12.32 2.40 12.32 1.54
                 0.51 1.54 0.51 1.22 17.78 1.22 17.78 1.54 12.64 1.54
                 12.64 2.08 13.06 2.08 13.06 3.58 14.14 3.58 14.14 2.94
                 14.46 2.94 14.46 3.58 15.54 3.58 15.54 2.94 15.86 2.94
                 15.86 3.58 16.94 3.58 16.94 2.94 17.26 2.94 17.26 3.58
                 18.34 3.58 18.34 2.94 18.66 2.94 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 19.20 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  19.20 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 3.58 1.20 3.58
                 1.20 4.86 2.28 4.86 2.28 3.58 2.60 3.58 2.60 4.86 3.68 4.86
                 3.68 3.58 4.00 3.58 4.00 4.86 5.08 4.86 5.08 4.22 5.40 4.22
                 5.40 4.86 19.20 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  17.98 4.54 12.06 4.54 12.06 3.90 6.46 3.90 6.46 2.94 6.78 2.94
                 6.78 3.58 7.86 3.58 7.86 2.94 8.18 2.94 8.18 3.58 9.26 3.58
                 9.26 2.94 9.58 2.94 9.58 3.58 10.66 3.58 10.66 2.94 10.98 2.94
                 10.98 3.58 12.06 3.58 12.06 2.94 12.38 2.94 12.38 4.22
                 17.98 4.22 ;
        POLYGON  11.69 4.54 5.78 4.54 5.78 3.90 4.70 3.90 4.70 4.54 4.38 4.54
                 4.38 3.26 3.30 3.26 3.30 4.54 2.98 4.54 2.98 3.26 1.90 3.26
                 1.90 4.54 1.58 4.54 1.58 3.26 0.50 3.26 0.50 4.54 0.18 4.54
                 0.18 2.94 4.70 2.94 4.70 3.58 6.10 3.58 6.10 4.22 11.69 4.22 ;
    END
END nor3_8

MACRO nor3_4
    CLASS CORE ;
    FOREIGN nor3_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.88 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  8.48 2.08 9.12 2.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.72 2.08 6.36 2.43 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.44 2.43 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 7.08  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.26 4.54 9.94 4.54 9.94 3.26 8.86 3.26 8.86 3.90 8.54 3.90
                 8.54 3.26 7.46 3.26 7.46 3.90 7.14 3.90 7.14 2.94 9.94 2.94
                 9.94 2.40 9.76 2.40 9.76 2.08 9.94 2.08 9.94 1.54 1.56 1.54
                 1.56 1.22 10.26 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 10.88 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  10.88 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 3.58 1.20 3.58
                 1.20 4.86 2.28 4.86 2.28 3.58 2.60 3.58 2.60 4.86 10.88 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  9.56 4.54 6.46 4.54 6.46 3.26 5.38 3.26 5.38 3.90 5.06 3.90
                 5.06 3.26 3.98 3.26 3.98 3.90 3.66 3.90 3.66 2.94 6.78 2.94
                 6.78 4.22 7.84 4.22 7.84 3.58 8.16 3.58 8.16 4.22 9.24 4.22
                 9.24 3.58 9.56 3.58 ;
        POLYGON  6.08 4.54 2.98 4.54 2.98 3.26 1.90 3.26 1.90 4.54 1.58 4.54
                 1.58 3.26 0.50 3.26 0.50 4.54 0.18 4.54 0.18 2.94 3.30 2.94
                 3.30 4.22 4.36 4.22 4.36 3.58 4.68 3.58 4.68 4.22 5.76 4.22
                 5.76 3.58 6.08 3.58 ;
    END
END nor3_4

MACRO nor3_2
    CLASS CORE ;
    FOREIGN nor3_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.32  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.08 4.96 2.72 ;
        END
    END a
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.32  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.48 2.08 1.12 2.43 ;
        END
    END c
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.32  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.16 2.08 3.80 2.43 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.40  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  6.06 4.54 5.74 4.54 5.74 3.90 4.34 3.90 4.34 3.58 5.74 3.58
                 5.74 2.40 5.28 2.40 5.28 2.08 5.74 2.08 5.74 1.54 0.85 1.54
                 0.85 1.22 6.06 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 6.40 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 3.58 1.20 3.58
                 1.20 4.86 6.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  5.36 4.54 3.66 4.54 3.66 3.26 2.58 3.26 2.58 3.90 2.26 3.90
                 2.26 2.94 3.98 2.94 3.98 4.22 5.36 4.22 ;
        POLYGON  3.28 4.54 1.58 4.54 1.58 3.26 0.50 3.26 0.50 4.54 0.18 4.54
                 0.18 2.94 1.90 2.94 1.90 4.22 2.96 4.22 2.96 3.58 3.28 3.58 ;
    END
END nor3_2

MACRO nor3_1
    CLASS CORE ;
    FOREIGN nor3_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.48 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.08 3.04 2.72 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.76 2.08 2.40 2.43 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.48 2.08 1.12 2.43 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.96 4.54 3.64 4.54 3.64 2.40 3.36 2.40 3.36 2.08 3.64 2.08
                 3.64 1.54 1.22 1.54 1.22 1.22 3.96 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  4.48 0.90 0.84 0.90 0.84 1.54 0.52 1.54 0.52 0.90 0.00 0.90
                 0.00 -0.90 4.48 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  4.48 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 3.58 1.20 3.58
                 1.20 4.86 4.48 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  2.26 3.58 3.26 4.54 ;
        POLYGON  1.88 4.54 1.56 4.54 1.56 3.26 0.50 3.26 0.50 4.54 0.18 4.54
                 0.18 2.94 1.56 2.94 1.56 2.78 1.88 2.78 ;
    END
END nor3_1

MACRO nor2a_8
    CLASS CORE ;
    FOREIGN nor2a_8 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.20 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.76 2.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 5.30  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  15.51 2.08 16.24 2.43 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 11.31  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  17.98 1.54 12.38 1.54 12.38 3.90 12.06 3.90 12.06 1.54
                 8.80 1.54 8.80 2.78 12.06 2.78 12.06 3.10 10.98 3.10
                 10.98 3.90 10.66 3.90 10.66 3.10 9.58 3.10 9.58 3.89 9.26 3.89
                 9.26 3.10 8.18 3.10 8.18 3.90 7.86 3.90 7.86 3.10 6.78 3.10
                 6.78 4.54 6.46 4.54 6.46 2.78 8.48 2.78 8.48 1.54 6.46 1.54
                 6.46 1.22 17.98 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 19.20 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  19.20 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 3.79 1.20 3.79
                 1.20 4.86 2.28 4.86 2.28 3.79 2.60 3.79 2.60 4.86 3.68 4.86
                 3.68 3.79 4.00 3.79 4.00 4.86 5.08 4.86 5.08 3.79 5.40 3.79
                 5.40 4.86 13.44 4.86 13.44 3.57 13.76 3.57 13.76 4.86
                 14.84 4.86 14.84 3.57 15.16 3.57 15.16 4.86 16.24 4.86
                 16.24 3.57 16.56 3.57 16.56 4.86 17.64 4.86 17.64 3.57
                 17.96 3.57 17.96 4.86 19.20 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  18.66 4.53 18.34 4.53 18.34 3.10 17.26 3.10 17.26 4.53
                 16.94 4.53 16.94 3.10 15.86 3.10 15.86 4.53 15.54 4.53
                 15.54 3.10 14.46 3.10 14.46 4.53 14.14 4.53 14.14 3.10
                 13.06 3.10 13.06 4.54 7.16 4.54 7.16 3.43 7.48 3.43 7.48 4.22
                 8.56 4.22 8.56 3.43 8.88 3.43 8.88 4.22 9.96 4.22 9.96 3.43
                 10.28 3.43 10.28 4.22 11.36 4.22 11.36 3.43 11.68 3.43
                 11.68 4.22 12.74 4.22 12.74 2.78 18.66 2.78 ;
        POLYGON  7.90 2.43 6.10 2.43 6.10 4.24 5.78 4.24 5.78 1.54 3.30 1.54
                 3.30 3.13 5.78 3.13 5.78 3.45 4.70 3.45 4.70 4.24 4.38 4.24
                 4.38 3.45 3.30 3.45 3.30 4.24 2.98 4.24 2.98 3.45 1.90 3.45
                 1.90 4.24 1.58 4.24 1.58 3.45 0.50 3.45 0.50 4.24 0.18 4.24
                 0.18 3.13 2.98 3.13 2.98 1.54 0.18 1.54 0.18 1.22 6.10 1.22
                 6.10 2.08 7.90 2.08 ;
    END
END nor2a_8

MACRO nor2a_4
    CLASS CORE ;
    FOREIGN nor2a_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.88 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.79  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.76 2.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  7.11 2.08 7.84 2.43 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.32  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.58 1.54 6.24 1.54 6.24 2.78 6.78 2.78 6.78 3.90 6.46 3.90
                 6.46 3.10 5.38 3.10 5.38 3.90 5.06 3.90 5.06 3.10 3.98 3.10
                 3.98 4.54 3.66 4.54 3.66 2.78 5.92 2.78 5.92 1.54 3.66 1.54
                 3.66 1.22 9.58 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 10.88 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  10.88 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 3.79 1.20 3.79
                 1.20 4.86 2.28 4.86 2.28 3.79 2.60 3.79 2.60 4.86 7.84 4.86
                 7.84 3.57 8.16 3.57 8.16 4.86 9.24 4.86 9.24 3.57 9.56 3.57
                 9.56 4.86 10.88 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  10.26 4.53 9.94 4.53 9.94 3.10 8.86 3.10 8.86 4.53 8.54 4.53
                 8.54 3.10 7.46 3.10 7.46 4.54 4.36 4.54 4.36 3.43 4.68 3.43
                 4.68 4.22 5.76 4.22 5.76 3.43 6.08 3.43 6.08 4.22 7.14 4.22
                 7.14 2.78 10.26 2.78 ;
        POLYGON  5.10 2.43 3.30 2.43 3.30 4.24 2.98 4.24 2.98 3.45 1.90 3.45
                 1.90 4.24 1.58 4.24 1.58 3.45 0.50 3.45 0.50 4.24 0.18 4.24
                 0.18 3.13 2.98 3.13 2.98 1.54 0.18 1.54 0.18 1.22 3.30 1.22
                 3.30 2.08 5.10 2.08 ;
    END
END nor2a_4

MACRO nor2a_2
    CLASS CORE ;
    FOREIGN nor2a_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.89  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.81 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.32  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.31 2.08 5.04 2.43 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.82  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  5.38 1.54 3.68 1.54 3.68 2.78 3.98 2.78 3.98 3.90 3.66 3.90
                 3.66 3.10 2.58 3.10 2.58 3.90 2.26 3.90 2.26 2.78 3.36 2.78
                 3.36 1.54 2.26 1.54 2.26 1.22 5.38 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 6.40 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 3.79 1.20 3.79
                 1.20 4.86 5.04 4.86 5.04 3.57 5.36 3.57 5.36 4.86 6.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  6.06 4.53 5.74 4.53 5.74 3.10 4.66 3.10 4.66 4.54 2.96 4.54
                 2.96 3.43 3.28 3.43 3.28 4.22 4.34 4.22 4.34 2.78 6.06 2.78 ;
        POLYGON  3.03 2.43 1.90 2.43 1.90 4.24 1.58 4.24 1.58 3.45 0.50 3.45
                 0.50 4.24 0.18 4.24 0.18 3.13 1.58 3.13 1.58 1.54 0.18 1.54
                 0.18 1.22 1.90 1.22 1.90 2.11 3.03 2.11 ;
    END
END nor2a_2

MACRO nor2a_1
    CLASS CORE ;
    FOREIGN nor2a_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.84 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.45  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 1.85 1.12 2.49 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 1.92 1.84 2.49 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.71  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.68 3.04 3.52 3.04 3.52 4.54 3.20 4.54 3.20 2.72 3.36 2.72
                 3.36 1.82 2.16 1.82 2.16 1.22 2.48 1.22 2.48 1.50 3.68 1.50 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  3.84 0.90 3.18 0.90 3.18 1.18 2.86 1.18 2.86 0.90 1.78 0.90
                 1.78 1.19 0.88 1.19 0.88 0.90 0.00 0.90 0.00 -0.90 3.84 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  3.84 6.66 0.00 6.66 0.00 4.86 0.99 4.86 0.99 4.28 1.31 4.28
                 1.31 4.86 3.84 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  2.88 3.13 0.48 3.13 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.81 2.56 2.81
                 2.56 2.17 2.88 2.17 ;
        RECT  1.82 3.45 2.82 4.54 ;
    END
END nor2a_1

MACRO nor2_8
    CLASS CORE ;
    FOREIGN nor2_8 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.80 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 5.30  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.56 2.08 11.48 2.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 5.30  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.08 1.76 2.43 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 11.31  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.38 3.90 6.46 3.90 6.46 3.26 5.92 3.26 5.92 1.54 0.51 1.54
                 0.51 1.22 12.04 1.22 12.04 1.54 6.24 1.54 6.24 2.94 6.78 2.94
                 6.78 3.58 7.86 3.58 7.86 2.94 8.18 2.94 8.18 3.58 9.26 3.58
                 9.26 2.94 9.58 2.94 9.58 3.58 10.66 3.58 10.66 2.94 10.98 2.94
                 10.98 3.58 12.06 3.58 12.06 2.94 12.38 2.94 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 12.80 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  12.80 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 3.58 1.20 3.58
                 1.20 4.86 2.28 4.86 2.28 3.58 2.60 3.58 2.60 4.86 3.68 4.86
                 3.68 3.58 4.00 3.58 4.00 4.86 5.08 4.86 5.08 4.22 5.40 4.22
                 5.40 4.86 12.80 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  11.69 4.54 5.78 4.54 5.78 3.90 4.70 3.90 4.70 4.54 4.38 4.54
                 4.38 3.26 3.30 3.26 3.30 4.54 2.98 4.54 2.98 3.26 1.90 3.26
                 1.90 4.54 1.58 4.54 1.58 3.26 0.50 3.26 0.50 4.54 0.18 4.54
                 0.18 2.94 4.70 2.94 4.70 3.58 6.10 3.58 6.10 4.22 11.69 4.22 ;
    END
END nor2_8

MACRO nor2_4
    CLASS CORE ;
    FOREIGN nor2_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.04 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.96 2.08 5.60 2.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.08 1.76 2.43 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.32  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  6.78 4.54 6.46 4.54 6.46 3.90 3.66 3.90 3.66 3.26 3.32 3.26
                 3.32 1.54 0.52 1.54 0.52 1.22 6.44 1.22 6.44 1.54 3.64 1.54
                 3.64 2.72 3.68 2.72 3.68 2.94 3.98 2.94 3.98 3.58 5.06 3.58
                 5.06 2.94 5.38 2.94 5.38 3.58 6.46 3.58 6.46 2.94 6.78 2.94 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 7.04 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.04 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 3.58 1.20 3.58
                 1.20 4.86 2.28 4.86 2.28 4.22 2.60 4.22 2.60 4.86 7.04 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  6.08 4.54 2.98 4.54 2.98 3.90 1.90 3.90 1.90 4.54 1.58 4.54
                 1.58 3.26 0.50 3.26 0.50 4.54 0.18 4.54 0.18 2.94 1.90 2.94
                 1.90 3.58 3.30 3.58 3.30 4.22 6.08 4.22 ;
    END
END nor2_4

MACRO nor2_2
    CLASS CORE ;
    FOREIGN nor2_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.48 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.32  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.04 2.08 3.68 2.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.32  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.08 1.76 2.43 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.83  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.22 4.54 3.90 4.54 3.90 3.90 2.50 3.90 2.50 3.26 2.16 3.26
                 2.16 3.04 2.08 3.04 2.08 2.72 2.16 2.72 2.16 1.54 0.76 1.54
                 0.76 1.22 3.88 1.22 3.88 1.54 2.48 1.54 2.48 2.94 2.82 2.94
                 2.82 3.58 3.90 3.58 3.90 2.94 4.22 2.94 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 4.48 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  4.48 6.66 0.00 6.66 0.00 4.86 0.42 4.86 0.42 3.58 0.74 3.58
                 0.74 4.86 4.48 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  3.52 4.54 1.12 4.54 1.12 2.94 1.44 2.94 1.44 4.22 3.52 4.22 ;
    END
END nor2_2

MACRO nor2_1
    CLASS CORE ;
    FOREIGN nor2_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.20 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.08 2.72 2.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.48 2.08 1.12 2.43 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.71  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  2.80 4.54 2.48 4.54 2.48 3.90 1.44 3.90 1.44 1.22 1.76 1.22
                 1.76 3.58 2.48 3.58 2.48 2.94 2.80 2.94 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  3.20 0.90 2.46 0.90 2.46 1.54 2.14 1.54 2.14 0.90 1.06 0.90
                 1.06 1.54 0.74 1.54 0.74 0.90 0.00 0.90 0.00 -0.90 3.20 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 3.20 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  2.10 4.54 0.40 4.54 0.40 2.94 0.72 2.94 0.72 4.22 2.10 4.22 ;
    END
END nor2_1

MACRO nand4_8
    CLASS CORE ;
    FOREIGN nand4_8 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.16 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.60 1.12 3.24 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.72 1.76 3.39 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.58  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.44 2.46 3.04 2.46 3.04 2.40 2.72 2.40 2.72 2.08 3.44 2.08 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.58  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.72 2.74 3.16 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.29  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  11.87 1.74 10.47 1.74 10.47 2.72 10.72 2.72 10.72 3.04
                 10.47 3.04 10.47 3.78 11.55 3.78 11.55 3.10 11.87 3.10
                 11.87 4.10 8.75 4.10 8.75 3.16 9.07 3.16 9.07 3.78 10.15 3.78
                 10.15 1.74 8.75 1.74 8.75 1.42 11.87 1.42 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  12.16 0.90 2.58 0.90 2.58 1.54 2.26 1.54 2.26 0.90 0.00 0.90
                 0.00 -0.90 12.16 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  12.16 6.66 0.00 6.66 0.00 4.86 9.45 4.86 9.45 4.42 9.77 4.42
                 9.77 4.86 10.85 4.86 10.85 4.42 11.17 4.42 11.17 4.86
                 12.16 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  9.69 2.66 8.39 2.66 8.39 4.54 8.07 4.54 8.07 3.90 6.67 3.90
                 6.67 3.58 8.07 3.58 8.07 1.54 5.03 1.54 5.03 1.22 8.39 1.22
                 8.39 2.34 9.69 2.34 ;
        POLYGON  7.69 4.54 5.29 4.54 5.29 3.58 5.61 3.58 5.61 4.22 7.69 4.22 ;
        POLYGON  7.09 3.25 4.83 3.25 4.83 3.90 4.31 3.90 4.31 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.56 0.48 1.56 0.48 4.22 3.99 4.22
                 3.99 3.58 4.51 3.58 4.51 2.93 6.77 2.93 6.77 2.11 7.09 2.11 ;
        POLYGON  5.93 2.43 4.08 2.43 4.08 3.10 3.52 3.10 3.52 3.90 3.20 3.90
                 3.20 2.78 3.76 2.78 3.76 2.08 4.34 2.08 4.34 1.22 4.66 1.22
                 4.66 2.11 5.93 2.11 ;
        RECT  2.96 1.22 3.96 1.54 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END nand4_8

MACRO nand4_4
    CLASS CORE ;
    FOREIGN nand4_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.96 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.60 1.12 3.24 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.72 1.76 3.39 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.58  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.44 2.46 3.04 2.46 3.04 2.40 2.72 2.40 2.72 2.08 3.44 2.08 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.58  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.72 2.74 3.16 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.77  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.62 4.54 8.30 4.54 8.30 3.68 7.22 3.68 7.22 4.54 6.90 4.54
                 6.90 3.36 8.30 3.36 8.30 1.70 7.35 1.70 7.35 1.38 8.62 1.38 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.96 0.90 2.58 0.90 2.58 1.54 2.26 1.54 2.26 0.90 0.00 0.90
                 0.00 -0.90 8.96 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  8.96 6.66 0.00 6.66 0.00 4.86 7.60 4.86 7.60 4.22 7.92 4.22
                 7.92 4.86 8.96 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  7.73 2.94 6.54 2.94 6.54 4.54 6.22 4.54 6.22 1.54 5.71 1.54
                 5.71 1.22 6.54 1.22 6.54 2.62 7.73 2.62 ;
        RECT  4.84 4.22 5.84 4.54 ;
        POLYGON  5.56 2.62 5.46 2.62 5.46 3.90 4.52 3.90 4.52 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.56 0.48 1.56 0.48 4.22 4.20 4.22
                 4.20 3.58 5.14 3.58 5.14 2.30 5.56 2.30 ;
        POLYGON  4.82 2.60 4.08 2.60 4.08 3.10 3.52 3.10 3.52 3.90 3.20 3.90
                 3.20 2.78 3.76 2.78 3.76 2.28 4.34 2.28 4.34 1.22 4.66 1.22
                 4.66 2.28 4.82 2.28 ;
        RECT  2.96 1.22 3.96 1.54 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END nand4_4

MACRO nand4_2
    CLASS CORE ;
    FOREIGN nand4_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.32 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.60 1.12 3.24 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.72 1.76 3.39 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.58  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.44 2.46 3.04 2.46 3.04 2.40 2.72 2.40 2.72 2.08 3.44 2.08 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.58  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.72 2.74 3.16 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.12 4.34 7.80 4.34 7.80 3.68 7.20 3.68 7.20 3.36 7.80 3.36
                 7.80 1.38 8.12 1.38 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 0.90 7.42 0.90 7.42 1.32 7.10 1.32 7.10 0.90 2.58 0.90
                 2.58 1.54 2.26 1.54 2.26 0.90 0.00 0.90 0.00 -0.90 8.32 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 8.32 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  7.10 2.94 6.54 2.94 6.54 4.54 6.22 4.54 6.22 1.54 5.02 1.54
                 5.02 1.22 6.74 1.22 6.74 1.54 6.54 1.54 6.54 2.62 7.10 2.62 ;
        RECT  4.84 4.22 5.84 4.54 ;
        POLYGON  5.56 2.62 5.46 2.62 5.46 3.90 4.52 3.90 4.52 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.56 0.48 1.56 0.48 4.22 4.20 4.22
                 4.20 3.58 5.14 3.58 5.14 2.30 5.56 2.30 ;
        POLYGON  4.82 2.60 4.08 2.60 4.08 3.10 3.52 3.10 3.52 3.90 3.20 3.90
                 3.20 2.78 3.76 2.78 3.76 2.28 4.34 2.28 4.34 1.22 4.66 1.22
                 4.66 2.28 4.82 2.28 ;
        RECT  2.96 1.22 3.96 1.54 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END nand4_2

MACRO nand4_1
    CLASS CORE ;
    FOREIGN nand4_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.32 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.60 1.12 3.24 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.72 1.76 3.39 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.58  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.44 2.46 3.04 2.46 3.04 2.40 2.72 2.40 2.72 2.08 3.44 2.08 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.58  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.72 2.74 3.16 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.12 4.34 7.80 4.34 7.80 3.68 7.20 3.68 7.20 3.36 7.80 3.36
                 7.80 1.38 8.12 1.38 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 0.90 7.42 0.90 7.42 1.32 7.10 1.32 7.10 0.90 2.58 0.90
                 2.58 1.54 2.26 1.54 2.26 0.90 0.00 0.90 0.00 -0.90 8.32 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 6.66 0.00 6.66 0.00 4.86 7.10 4.86 7.10 4.34 7.42 4.34
                 7.42 4.86 8.32 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  7.10 2.94 6.54 2.94 6.54 4.54 6.22 4.54 6.22 1.54 5.02 1.54
                 5.02 1.22 6.74 1.22 6.74 1.54 6.54 1.54 6.54 2.62 7.10 2.62 ;
        RECT  4.84 4.22 5.84 4.54 ;
        POLYGON  5.56 2.62 5.46 2.62 5.46 3.90 4.52 3.90 4.52 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.56 0.48 1.56 0.48 4.22 4.20 4.22
                 4.20 3.58 5.14 3.58 5.14 2.30 5.56 2.30 ;
        POLYGON  4.82 2.60 4.08 2.60 4.08 3.10 3.52 3.10 3.52 3.90 3.20 3.90
                 3.20 2.78 3.76 2.78 3.76 2.28 4.34 2.28 4.34 1.22 4.66 1.22
                 4.66 2.28 4.82 2.28 ;
        RECT  2.96 1.22 3.96 1.54 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END nand4_1

MACRO nand3_8
    CLASS CORE ;
    FOREIGN nand3_8 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.20 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 4.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 2.62 5.60 3.26 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 4.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.48 2.62 6.98 3.26 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 4.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  12.96 2.72 13.56 3.26 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 14.48  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  17.75 4.54 4.64 4.54 4.64 2.22 1.12 2.22 1.12 4.22 4.64 4.22
                 4.64 4.54 0.52 4.54 0.52 4.22 0.80 4.22 0.80 2.22 0.18 2.22
                 0.18 1.90 6.10 1.90 6.10 2.22 4.96 2.22 4.96 4.22 17.75 4.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 19.20 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 19.20 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  18.70 1.92 13.06 1.92 13.06 2.22 7.16 2.22 7.16 1.90
                 12.74 1.90 12.74 1.60 18.70 1.60 ;
        RECT  0.87 1.22 12.38 1.54 ;
    END
END nand3_8

MACRO nand3_4
    CLASS CORE ;
    FOREIGN nand3_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.88 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.26  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.18 2.72 1.76 3.37 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.26  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.72 4.96 3.37 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.26  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  8.48 2.72 8.80 3.37 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 8.88  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.26 4.54 0.18 4.54 0.18 1.22 0.50 1.22 0.50 1.86 3.30 1.86
                 3.30 2.18 0.50 2.18 0.50 4.22 9.12 4.22 9.12 4.00 9.44 4.00
                 9.44 4.22 10.26 4.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 10.88 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 10.88 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  4.36 1.22 10.26 1.54 ;
        POLYGON  6.78 2.18 3.62 2.18 3.62 1.54 0.88 1.54 0.88 1.22 3.94 1.22
                 3.94 1.86 6.78 1.86 ;
    END
END nand3_4

MACRO nand3_2
    CLASS CORE ;
    FOREIGN nand3_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.13  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.18 2.72 1.76 3.37 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.13  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.04 3.37 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.13  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.72 4.96 3.37 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.58  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  6.06 4.54 0.18 4.54 0.18 1.22 0.50 1.22 0.50 1.86 1.90 1.86
                 1.90 2.18 0.50 2.18 0.50 4.22 5.28 4.22 5.28 4.00 5.60 4.00
                 5.60 4.22 6.06 4.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 6.40 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 6.40 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  2.96 1.22 6.06 1.54 ;
        POLYGON  3.98 2.18 2.26 2.18 2.26 1.54 0.88 1.54 0.88 1.22 2.58 1.22
                 2.58 1.86 3.98 1.86 ;
    END
END nand3_2

MACRO nand3_1
    CLASS CORE ;
    FOREIGN nand3_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.48 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.62 1.12 3.26 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.62 1.76 3.26 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.04 3.37 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.21  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.04 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.56 0.48 1.56
                 0.48 4.22 3.04 4.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  4.48 0.90 3.96 0.90 3.96 1.54 3.64 1.54 3.64 0.90 0.00 0.90
                 0.00 -0.90 4.48 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 4.48 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  2.26 1.22 3.26 1.54 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END nand3_1

MACRO nand2a_8
    CLASS CORE ;
    FOREIGN nand2a_8 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.64 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.79  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.72 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 4.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  13.06 2.72 13.96 3.04 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 10.99  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  15.26 4.36 3.65 4.36 3.65 4.04 9.12 4.04 9.12 2.18 3.66 2.18
                 3.66 1.86 9.58 1.86 9.58 2.18 9.44 2.18 9.44 4.04 15.26 4.04 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 16.88 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.88 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 3.91 1.20 3.91
                 1.20 4.86 2.27 4.86 2.27 3.90 2.60 3.90 2.60 4.86 4.36 4.86
                 4.36 4.68 4.68 4.68 4.68 4.86 5.76 4.86 5.76 4.68 6.08 4.68
                 6.08 4.86 7.16 4.86 7.16 4.68 7.48 4.68 7.48 4.86 8.56 4.86
                 8.56 4.68 8.89 4.68 8.89 4.86 9.97 4.86 9.97 4.68 10.29 4.68
                 10.29 4.86 11.39 4.86 11.39 4.68 11.72 4.68 11.72 4.86
                 12.81 4.86 12.81 4.68 13.14 4.68 13.14 4.86 14.23 4.86
                 14.23 4.68 14.56 4.68 14.56 4.86 16.88 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  4.35 1.22 15.94 1.54 ;
        POLYGON  5.03 3.58 2.97 3.58 2.97 1.54 1.89 1.54 1.89 3.26 2.97 3.26
                 2.97 3.58 0.16 3.58 0.16 3.26 1.56 3.26 1.56 1.54 0.16 1.54
                 0.16 1.22 3.30 1.22 3.30 3.26 5.03 3.26 ;
    END
END nand2a_8

MACRO nand2a_4
    CLASS CORE ;
    FOREIGN nand2a_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.60 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.89  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.72 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.26  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  7.08 2.72 7.72 3.04 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.06  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.22 4.36 2.24 4.36 2.24 4.04 4.64 4.04 4.64 2.18 2.26 2.18
                 2.26 1.86 5.38 1.86 5.38 2.18 4.96 2.18 4.96 4.04 8.22 4.04 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 9.60 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  9.60 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 3.91 1.20 3.91
                 1.20 4.86 2.96 4.86 2.96 4.68 3.28 4.68 3.28 4.86 4.36 4.86
                 4.36 4.68 4.69 4.68 4.69 4.86 5.77 4.86 5.77 4.68 6.09 4.68
                 6.09 4.86 7.19 4.86 7.19 4.68 7.52 4.68 7.52 4.86 9.60 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  2.95 1.22 8.90 1.54 ;
        POLYGON  2.67 3.58 0.16 3.58 0.16 3.26 1.57 3.26 1.57 1.54 0.16 1.54
                 0.16 1.22 1.90 1.22 1.90 3.26 2.67 3.26 ;
    END
END nand2a_4

MACRO nand2a_2
    CLASS CORE ;
    FOREIGN nand2a_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.89  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.72 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.13  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.48 2.72 5.12 3.04 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.17  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  6.08 4.36 2.24 4.36 2.24 4.04 3.36 4.04 3.36 2.83 2.24 2.83
                 2.24 1.22 3.98 1.22 3.98 1.54 2.56 1.54 2.56 2.51 3.68 2.51
                 3.68 4.04 6.08 4.04 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 0.90 5.37 0.90 5.37 1.08 5.05 1.08 5.05 0.90 1.20 0.90
                 1.20 1.66 0.88 1.66 0.88 0.90 0.00 0.90 0.00 -0.90 6.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.66 1.20 4.66
                 1.20 4.86 2.96 4.86 2.96 4.68 3.28 4.68 3.28 4.86 5.05 4.86
                 5.05 4.68 5.37 4.68 5.37 4.86 6.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  6.08 1.72 4.62 1.72 4.62 2.18 2.96 2.18 2.96 1.86 4.30 1.86
                 4.30 1.40 6.08 1.40 ;
        POLYGON  2.48 3.58 1.92 3.58 1.92 4.54 1.58 4.54 1.58 4.22 1.60 4.22
                 1.60 3.58 0.48 3.58 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 3.26 1.60 3.26
                 1.60 1.54 1.58 1.54 1.58 1.22 1.92 1.22 1.92 3.26 2.48 3.26 ;
    END
END nand2a_2

MACRO nand2a_1
    CLASS CORE ;
    FOREIGN nand2a_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.84 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.45  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.04 3.04 2.68 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.04 2.40 2.68 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.98 4.36 0.28 4.36 0.28 3.72 0.16 3.72 0.16 2.10 0.28 2.10
                 0.28 1.22 0.60 1.22 0.60 2.42 0.48 2.42 0.48 3.40 0.60 3.40
                 0.60 4.04 1.98 4.04 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 3.84 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 3.84 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  3.68 4.36 3.30 4.36 3.30 4.04 3.36 4.04 3.36 3.58 0.92 3.58
                 0.92 3.26 3.36 3.26 3.36 1.54 3.30 1.54 3.30 1.22 3.68 1.22 ;
        RECT  0.98 1.22 1.98 1.54 ;
    END
END nand2a_1

MACRO nand2_8
    CLASS CORE ;
    FOREIGN nand2_8 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.80 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 4.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 2.62 5.60 3.26 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 4.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.48 2.62 6.98 3.26 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 10.99  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.04 4.54 4.64 4.54 4.64 2.22 1.12 2.22 1.12 4.22 4.64 4.22
                 4.64 4.54 0.52 4.54 0.52 4.22 0.80 4.22 0.80 2.22 0.18 2.22
                 0.18 1.90 6.10 1.90 6.10 2.22 4.96 2.22 4.96 4.22 12.04 4.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 12.80 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 12.80 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  0.87 1.22 12.38 1.54 ;
    END
END nand2_8

MACRO nand2_4
    CLASS CORE ;
    FOREIGN nand2_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.04 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.26  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.62 3.04 3.26 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.26  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.62 3.86 3.26 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.06  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  6.44 4.54 0.52 4.54 0.52 4.22 2.08 4.22 2.08 2.22 0.18 2.22
                 0.18 1.22 0.50 1.22 0.50 1.90 3.30 1.90 3.30 2.22 2.40 2.22
                 2.40 4.22 6.44 4.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 7.04 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 7.04 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  0.88 1.22 6.78 1.54 ;
    END
END nand2_4

MACRO nand2_2
    CLASS CORE ;
    FOREIGN nand2_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.48 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.13  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.62 1.76 3.26 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.13  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.62 2.46 3.26 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.64 4.54 0.52 4.54 0.52 4.22 0.80 4.22 0.80 2.22 0.18 2.22
                 0.18 1.22 0.50 1.22 0.50 1.90 1.90 1.90 1.90 2.22 1.12 2.22
                 1.12 4.22 3.64 4.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 4.48 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 4.48 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  0.88 1.22 3.98 1.54 ;
    END
END nand2_2

MACRO nand2_1
    CLASS CORE ;
    FOREIGN nand2_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.20 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.62 1.12 3.26 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.62 1.76 3.26 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.51  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.44 4.54 1.12 4.54 1.12 3.90 0.16 3.90 0.16 1.22 0.50 1.22
                 0.50 1.56 0.48 1.56 0.48 3.58 1.44 3.58 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  3.20 0.90 2.58 0.90 2.58 1.54 2.26 1.54 2.26 0.90 0.00 0.90
                 0.00 -0.90 3.20 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  3.20 6.66 0.00 6.66 0.00 4.86 0.42 4.86 0.42 4.22 0.74 4.22
                 0.74 4.86 1.82 4.86 1.82 4.22 2.14 4.22 2.14 4.86 3.20 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END nand2_1

MACRO muxi8_4
    CLASS CORE ;
    FOREIGN muxi8_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 41.60 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.62 2.52 3.26 ;
        END
    END d0
    PIN d1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.96 2.72 3.68 3.12 ;
        END
    END d1
    PIN d2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.40 2.72 10.94 3.16 ;
        END
    END d2
    PIN d3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  9.12 2.54 9.44 3.18 ;
        END
    END d3
    PIN d4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  27.04 2.62 27.55 3.06 ;
        END
    END d4
    PIN d5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  26.24 2.62 26.72 3.06 ;
        END
    END d5
    PIN d6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  18.72 2.62 19.16 3.26 ;
        END
    END d6
    PIN d7
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  19.62 2.72 20.32 3.26 ;
        END
    END d7
    PIN sl0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.56 3.04 13.68 3.04 13.68 2.47 14.00 2.47 14.00 2.72
                 14.56 2.72 ;
        END
    END sl0
    PIN sl1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.98  LAYER metal1  ;
        ANTENNAGATEAREA 2.11  LAYER metal2  ;
        ANTENNAMAXAREACAR 0.02  LAYER metal1  ;
        ANTENNAMAXAREACAR 0.39  LAYER metal2  ;
        PORT
        LAYER metal2 ;
                POLYGON  22.36 3.90 6.76 3.90 6.76 2.74 7.08 2.74 7.08 3.58 15.76 3.58
                 15.76 2.72 16.08 2.72 16.08 3.58 22.04 3.58 22.04 2.72
                 22.36 2.72 ;
        LAYER v1 ;
        RECT  22.04 2.72 22.36 3.04 ;
        RECT  15.76 2.72 16.08 3.04 ;
        RECT  6.76 2.74 7.08 3.06 ;
        LAYER metal1 ;
        RECT  22.04 2.35 22.36 3.04 ;
        RECT  15.52 2.62 16.08 3.26 ;
        RECT  6.76 2.37 7.08 3.06 ;
        END
    END sl1
    PIN sl2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.18  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  31.96 3.68 31.52 3.68 31.52 3.36 31.64 3.36 31.64 2.62
                 31.96 2.62 ;
        END
    END sl2
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  41.42 4.32 39.70 4.32 39.70 4.00 41.10 4.00 41.10 1.59
                 39.70 1.59 39.70 1.27 41.42 1.27 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  41.60 0.90 26.94 0.90 26.94 1.14 26.62 1.14 26.62 0.90
                 19.54 0.90 19.54 1.14 19.22 1.14 19.22 0.90 16.08 0.90
                 16.08 1.14 15.76 1.14 15.76 0.90 14.00 0.90 14.00 1.14
                 13.68 1.14 13.68 0.90 10.54 0.90 10.54 1.14 10.22 1.14
                 10.22 0.90 2.98 0.90 2.98 1.14 2.66 1.14 2.66 0.90 0.00 0.90
                 0.00 -0.90 41.60 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  41.60 6.66 0.00 6.66 0.00 4.86 13.68 4.86 13.68 4.62
                 14.00 4.62 14.00 4.86 15.76 4.86 15.76 4.62 16.08 4.62
                 16.08 4.86 41.60 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  40.68 2.68 39.34 2.68 39.34 3.92 39.02 3.92 39.02 1.63
                 39.34 1.63 39.34 2.36 40.68 2.36 ;
        RECT  38.38 1.44 38.70 2.45 ;
        POLYGON  37.96 4.39 37.64 4.39 37.64 3.08 36.30 3.08 36.30 2.36
                 36.62 2.36 36.62 2.76 37.64 2.76 37.64 1.22 37.96 1.22 ;
        RECT  37.00 1.77 37.32 2.44 ;
        RECT  35.32 1.22 36.32 1.54 ;
        RECT  35.32 4.14 36.32 4.46 ;
        POLYGON  35.10 3.82 34.94 3.82 34.94 4.54 32.56 4.54 32.56 4.22
                 34.62 4.22 34.62 3.50 34.78 3.50 34.78 2.18 34.62 2.18
                 34.62 1.44 34.94 1.44 34.94 1.86 35.10 1.86 ;
        POLYGON  34.46 3.04 33.56 3.04 33.56 3.90 33.24 3.90 33.24 2.44
                 32.26 2.44 32.26 2.12 33.24 2.12 33.24 1.22 33.56 1.22
                 33.56 2.72 34.46 2.72 ;
        RECT  32.50 1.22 32.88 1.80 ;
        RECT  31.18 1.22 32.18 1.54 ;
        RECT  31.18 4.14 32.18 4.46 ;
        POLYGON  31.10 3.08 29.86 3.08 29.86 4.06 29.54 4.06 29.54 1.22
                 29.86 1.22 29.86 2.76 30.78 2.76 30.78 2.62 31.10 2.62 ;
        RECT  30.18 1.54 30.50 2.44 ;
        RECT  21.98 4.22 29.18 4.54 ;
        POLYGON  29.02 2.18 24.54 2.18 24.54 1.78 23.38 1.78 23.38 1.46
                 24.86 1.46 24.86 1.86 28.70 1.86 28.70 1.46 29.02 1.46 ;
        RECT  27.46 3.38 28.48 3.70 ;
        RECT  28.00 2.50 28.46 3.06 ;
        RECT  27.32 1.22 28.32 1.54 ;
        RECT  25.40 3.38 26.40 3.70 ;
        RECT  25.24 1.22 26.24 1.54 ;
        RECT  25.25 2.64 25.78 3.06 ;
        RECT  24.18 2.98 24.50 3.68 ;
        RECT  17.14 3.58 23.86 3.90 ;
        POLYGON  23.08 3.25 22.68 3.25 22.68 1.58 23.00 1.58 23.00 2.93
                 23.08 2.93 ;
        POLYGON  22.30 1.78 21.62 1.78 21.62 2.18 17.14 2.18 17.14 1.46
                 17.46 1.46 17.46 1.86 21.30 1.86 21.30 1.46 22.30 1.46 ;
        RECT  20.90 2.62 21.22 3.26 ;
        RECT  19.92 1.22 20.92 1.54 ;
        RECT  19.92 4.22 20.92 4.54 ;
        RECT  17.84 1.22 18.84 1.54 ;
        RECT  17.82 4.22 18.84 4.54 ;
        RECT  18.00 2.62 18.32 3.26 ;
        POLYGON  16.79 4.54 16.47 4.54 16.47 4.30 15.38 4.30 15.38 4.54
                 15.06 4.54 15.06 3.98 16.47 3.98 16.47 1.90 15.06 1.90
                 15.06 1.58 16.79 1.58 ;
        POLYGON  14.70 1.90 13.30 1.90 13.30 3.38 14.70 3.38 14.70 3.70
                 12.98 3.70 12.98 1.44 13.30 1.44 13.30 1.58 14.70 1.58 ;
        POLYGON  12.62 2.18 7.50 2.18 7.50 1.78 6.82 1.78 6.82 1.46 7.82 1.46
                 7.82 1.86 12.30 1.86 12.30 1.46 12.62 1.46 ;
        POLYGON  12.62 3.90 7.82 3.90 7.82 4.54 5.25 4.54 5.25 4.22 7.50 4.22
                 7.50 3.58 12.62 3.58 ;
        RECT  10.92 4.22 11.94 4.54 ;
        RECT  10.92 1.22 11.92 1.54 ;
        RECT  11.44 2.61 11.76 3.26 ;
        RECT  8.20 1.22 9.84 1.54 ;
        RECT  8.20 4.22 9.84 4.54 ;
        RECT  7.80 2.50 8.12 3.14 ;
        POLYGON  7.14 3.90 0.42 3.90 0.42 3.58 6.82 3.58 6.82 3.38 7.14 3.38 ;
        POLYGON  6.44 3.26 6.12 3.26 6.12 3.25 6.04 3.25 6.04 2.93 6.12 2.93
                 6.12 1.22 6.44 1.22 ;
        POLYGON  5.74 1.78 5.06 1.78 5.06 2.18 0.58 2.18 0.58 1.46 0.90 1.46
                 0.90 1.86 4.74 1.86 4.74 1.46 5.74 1.46 ;
        RECT  5.08 2.90 5.72 3.22 ;
        RECT  4.15 2.64 4.50 3.25 ;
        RECT  3.36 1.22 4.36 1.54 ;
        RECT  3.20 4.22 4.20 4.54 ;
        RECT  1.28 1.22 2.28 1.54 ;
        RECT  1.12 4.22 2.14 4.54 ;
        RECT  1.28 2.50 1.60 3.14 ;
        LAYER v1 ;
        RECT  38.38 1.44 38.70 1.76 ;
        RECT  37.00 2.12 37.32 2.44 ;
        RECT  34.62 1.44 34.94 1.76 ;
        RECT  32.56 1.44 32.88 1.76 ;
        RECT  30.18 1.54 30.50 1.86 ;
        RECT  28.00 2.50 28.32 2.82 ;
        RECT  25.46 2.64 25.78 2.96 ;
        RECT  24.18 3.36 24.50 3.68 ;
        RECT  22.68 2.72 23.00 3.04 ;
        RECT  20.90 2.64 21.22 2.96 ;
        RECT  18.00 2.64 18.32 2.96 ;
        RECT  16.47 4.22 16.79 4.54 ;
        RECT  15.06 4.22 15.38 4.54 ;
        RECT  12.98 1.86 13.30 2.18 ;
        RECT  11.44 2.66 11.76 2.98 ;
        RECT  7.80 2.66 8.12 2.98 ;
        RECT  6.12 1.22 6.44 1.54 ;
        RECT  5.40 2.90 5.72 3.22 ;
        RECT  4.18 2.64 4.50 2.96 ;
        RECT  1.28 2.50 1.60 2.82 ;
        LAYER metal2 ;
        RECT  32.56 1.44 38.70 1.76 ;
        POLYGON  37.32 4.32 24.82 4.32 24.82 3.04 22.68 3.04 22.68 2.72
                 25.14 2.72 25.14 4.00 37.00 4.00 37.00 2.12 37.32 2.12 ;
        POLYGON  30.50 1.86 30.18 1.86 30.18 1.54 6.12 1.54 6.12 1.22
                 30.50 1.22 ;
        POLYGON  28.32 2.82 28.00 2.82 28.00 2.18 25.78 2.18 25.78 2.96
                 25.46 2.96 25.46 2.18 21.22 2.18 21.22 2.96 20.90 2.96
                 20.90 2.18 18.32 2.18 18.32 2.96 18.00 2.96 18.00 2.18
                 11.76 2.18 11.76 2.98 11.44 2.98 11.44 2.18 8.12 2.18
                 8.12 2.98 7.80 2.98 7.80 2.18 4.50 2.18 4.50 2.96 4.18 2.96
                 4.18 2.18 1.60 2.18 1.60 2.82 1.28 2.82 1.28 1.86 28.32 1.86 ;
        POLYGON  24.50 4.54 5.40 4.54 5.40 2.90 5.72 2.90 5.72 4.22 24.18 4.22
                 24.18 3.36 24.50 3.36 ;
    END
END muxi8_4

MACRO muxi8_2
    CLASS CORE ;
    FOREIGN muxi8_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 40.96 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.62 2.52 3.26 ;
        END
    END d0
    PIN d1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.96 2.72 3.68 3.12 ;
        END
    END d1
    PIN d2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.40 2.72 10.94 3.16 ;
        END
    END d2
    PIN d3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  9.12 2.54 9.44 3.18 ;
        END
    END d3
    PIN d4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  27.04 2.62 27.46 3.26 ;
        END
    END d4
    PIN d5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  26.30 2.62 26.72 3.26 ;
        END
    END d5
    PIN d6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  18.72 2.62 19.16 3.26 ;
        END
    END d6
    PIN d7
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  19.62 2.72 20.32 3.26 ;
        END
    END d7
    PIN sl0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.56 3.04 13.68 3.04 13.68 2.47 14.00 2.47 14.00 2.72
                 14.56 2.72 ;
        END
    END sl0
    PIN sl1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.98  LAYER metal1  ;
        ANTENNAGATEAREA 2.11  LAYER metal2  ;
        ANTENNAMAXAREACAR 0.02  LAYER metal1  ;
        ANTENNAMAXAREACAR 0.39  LAYER metal2  ;
        PORT
        LAYER metal2 ;
                POLYGON  22.36 3.90 6.76 3.90 6.76 2.74 7.08 2.74 7.08 3.58 15.76 3.58
                 15.76 2.72 16.08 2.72 16.08 3.58 22.04 3.58 22.04 2.72
                 22.36 2.72 ;
        LAYER v1 ;
        RECT  22.04 2.72 22.36 3.04 ;
        RECT  15.76 2.72 16.08 3.04 ;
        RECT  6.76 2.74 7.08 3.06 ;
        LAYER metal1 ;
        RECT  22.04 2.35 22.36 3.04 ;
        RECT  15.52 2.62 16.08 3.26 ;
        RECT  6.76 2.37 7.08 3.06 ;
        END
    END sl1
    PIN sl2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.18  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  32.02 3.68 31.52 3.68 31.52 3.36 31.70 3.36 31.70 2.62
                 32.02 2.62 ;
        END
    END sl2
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  40.80 3.76 40.46 3.76 40.46 3.44 40.48 3.44 40.48 1.59
                 40.46 1.59 40.46 1.27 40.80 1.27 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  40.96 0.90 27.00 0.90 27.00 1.14 26.68 1.14 26.68 0.90
                 19.54 0.90 19.54 1.14 19.22 1.14 19.22 0.90 16.08 0.90
                 16.08 1.14 15.76 1.14 15.76 0.90 14.00 0.90 14.00 1.14
                 13.68 1.14 13.68 0.90 10.54 0.90 10.54 1.14 10.22 1.14
                 10.22 0.90 2.98 0.90 2.98 1.14 2.66 1.14 2.66 0.90 0.00 0.90
                 0.00 -0.90 40.96 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  40.96 6.66 0.00 6.66 0.00 4.86 13.68 4.86 13.68 4.62
                 14.00 4.62 14.00 4.86 15.76 4.86 15.76 4.62 16.08 4.62
                 16.08 4.86 40.96 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  40.16 2.68 39.40 2.68 39.40 3.92 39.08 3.92 39.08 1.63
                 39.40 1.63 39.40 2.36 40.16 2.36 ;
        RECT  38.44 1.44 38.76 2.45 ;
        POLYGON  38.02 4.39 37.70 4.39 37.70 3.08 36.46 3.08 36.46 2.62
                 36.78 2.62 36.78 2.76 37.70 2.76 37.70 1.22 38.02 1.22 ;
        RECT  37.06 1.80 37.38 2.44 ;
        RECT  35.38 1.22 36.38 1.54 ;
        RECT  35.38 4.14 36.38 4.46 ;
        POLYGON  35.16 3.82 35.00 3.82 35.00 4.54 32.62 4.54 32.62 4.22
                 34.68 4.22 34.68 3.50 34.84 3.50 34.84 2.18 34.68 2.18
                 34.68 1.36 35.00 1.36 35.00 1.86 35.16 1.86 ;
        POLYGON  34.52 3.04 33.62 3.04 33.62 3.90 33.30 3.90 33.30 2.44
                 32.32 2.44 32.32 2.12 33.30 2.12 33.30 1.22 33.62 1.22
                 33.62 2.72 34.52 2.72 ;
        RECT  32.56 1.22 32.94 1.80 ;
        RECT  31.24 1.22 32.24 1.54 ;
        RECT  31.24 4.14 32.24 4.46 ;
        POLYGON  31.16 3.08 29.92 3.08 29.92 4.06 29.60 4.06 29.60 1.22
                 29.92 1.22 29.92 2.76 30.84 2.76 30.84 2.62 31.16 2.62 ;
        RECT  30.24 1.22 30.56 2.44 ;
        POLYGON  29.24 3.90 25.14 3.90 25.14 4.54 21.98 4.54 21.98 4.22
                 24.82 4.22 24.82 3.58 29.24 3.58 ;
        POLYGON  29.08 2.18 24.60 2.18 24.60 1.78 23.38 1.78 23.38 1.46
                 24.92 1.46 24.92 1.86 28.76 1.86 28.76 1.46 29.08 1.46 ;
        RECT  27.52 4.22 28.54 4.54 ;
        RECT  27.38 1.22 28.38 1.54 ;
        RECT  28.06 2.50 28.38 3.14 ;
        RECT  25.46 4.22 26.46 4.54 ;
        RECT  25.30 1.22 26.30 1.54 ;
        RECT  25.46 2.62 25.78 3.26 ;
        RECT  24.18 3.24 24.50 3.90 ;
        RECT  17.14 3.58 23.86 3.90 ;
        POLYGON  23.08 3.25 22.68 3.25 22.68 1.58 23.00 1.58 23.00 2.93
                 23.08 2.93 ;
        POLYGON  22.30 1.78 21.62 1.78 21.62 2.18 17.14 2.18 17.14 1.46
                 17.46 1.46 17.46 1.86 21.30 1.86 21.30 1.46 22.30 1.46 ;
        RECT  20.90 2.62 21.22 3.26 ;
        RECT  19.92 1.22 20.92 1.54 ;
        RECT  19.92 4.22 20.92 4.54 ;
        RECT  17.84 1.22 18.84 1.54 ;
        RECT  17.82 4.22 18.84 4.54 ;
        RECT  18.00 2.62 18.32 3.26 ;
        POLYGON  16.79 4.54 16.47 4.54 16.47 4.30 15.38 4.30 15.38 4.54
                 15.06 4.54 15.06 3.98 16.47 3.98 16.47 1.90 15.06 1.90
                 15.06 1.58 16.79 1.58 ;
        POLYGON  14.70 1.90 13.30 1.90 13.30 3.38 14.70 3.38 14.70 3.70
                 12.98 3.70 12.98 1.44 13.30 1.44 13.30 1.58 14.70 1.58 ;
        POLYGON  12.62 2.18 7.50 2.18 7.50 1.78 6.82 1.78 6.82 1.46 7.82 1.46
                 7.82 1.86 12.30 1.86 12.30 1.46 12.62 1.46 ;
        POLYGON  12.62 3.90 7.82 3.90 7.82 4.54 5.25 4.54 5.25 4.22 7.50 4.22
                 7.50 3.58 12.62 3.58 ;
        RECT  10.92 4.22 11.94 4.54 ;
        RECT  10.92 1.22 11.92 1.54 ;
        RECT  11.44 2.61 11.76 3.26 ;
        RECT  8.20 1.22 9.84 1.54 ;
        RECT  8.20 4.22 9.84 4.54 ;
        RECT  7.80 2.50 8.12 3.14 ;
        POLYGON  7.14 3.90 0.42 3.90 0.42 3.58 6.82 3.58 6.82 3.38 7.14 3.38 ;
        POLYGON  6.44 3.26 6.12 3.26 6.12 3.25 6.04 3.25 6.04 2.93 6.12 2.93
                 6.12 1.22 6.44 1.22 ;
        POLYGON  5.74 1.78 5.06 1.78 5.06 2.18 0.58 2.18 0.58 1.46 0.90 1.46
                 0.90 1.86 4.74 1.86 4.74 1.46 5.74 1.46 ;
        RECT  5.08 2.90 5.72 3.22 ;
        RECT  4.15 2.64 4.50 3.25 ;
        RECT  3.36 1.22 4.36 1.54 ;
        RECT  3.20 4.22 4.20 4.54 ;
        RECT  1.28 1.22 2.28 1.54 ;
        RECT  1.12 4.22 2.14 4.54 ;
        RECT  1.28 2.50 1.60 3.14 ;
        LAYER v1 ;
        RECT  38.44 1.44 38.76 1.76 ;
        RECT  37.06 2.12 37.38 2.44 ;
        RECT  34.68 1.44 35.00 1.76 ;
        RECT  32.62 1.44 32.94 1.76 ;
        RECT  30.24 1.22 30.56 1.54 ;
        RECT  28.06 2.50 28.38 2.82 ;
        RECT  25.46 2.64 25.78 2.96 ;
        RECT  24.18 3.58 24.50 3.90 ;
        RECT  22.68 2.72 23.00 3.04 ;
        RECT  20.90 2.64 21.22 2.96 ;
        RECT  18.00 2.64 18.32 2.96 ;
        RECT  16.47 4.22 16.79 4.54 ;
        RECT  15.06 4.22 15.38 4.54 ;
        RECT  12.98 1.86 13.30 2.18 ;
        RECT  11.44 2.66 11.76 2.98 ;
        RECT  7.80 2.66 8.12 2.98 ;
        RECT  6.12 1.22 6.44 1.54 ;
        RECT  5.40 2.90 5.72 3.22 ;
        RECT  4.18 2.64 4.50 2.96 ;
        RECT  1.28 2.50 1.60 2.82 ;
        LAYER metal2 ;
        RECT  32.62 1.44 38.76 1.76 ;
        POLYGON  37.38 4.54 24.82 4.54 24.82 3.04 22.68 3.04 22.68 2.72
                 25.14 2.72 25.14 4.00 37.06 4.00 37.06 2.12 37.38 2.12 ;
        RECT  6.12 1.22 30.56 1.54 ;
        POLYGON  28.38 2.82 28.06 2.82 28.06 2.18 25.78 2.18 25.78 2.96
                 25.46 2.96 25.46 2.18 21.22 2.18 21.22 2.96 20.90 2.96
                 20.90 2.18 18.32 2.18 18.32 2.96 18.00 2.96 18.00 2.18
                 11.76 2.18 11.76 2.98 11.44 2.98 11.44 2.18 8.12 2.18
                 8.12 2.98 7.80 2.98 7.80 2.18 4.50 2.18 4.50 2.96 4.18 2.96
                 4.18 2.18 1.60 2.18 1.60 2.82 1.28 2.82 1.28 1.86 28.38 1.86 ;
        POLYGON  24.50 4.54 5.40 4.54 5.40 2.90 5.72 2.90 5.72 4.22 24.18 4.22
                 24.18 3.53 24.50 3.53 ;
    END
END muxi8_2

MACRO muxi8_1
    CLASS CORE ;
    FOREIGN muxi8_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 40.96 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.62 2.52 3.26 ;
        END
    END d0
    PIN d1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.96 2.72 3.68 3.12 ;
        END
    END d1
    PIN d2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.40 2.72 10.94 3.16 ;
        END
    END d2
    PIN d3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  9.12 2.54 9.44 3.18 ;
        END
    END d3
    PIN d4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  27.04 2.62 27.46 3.26 ;
        END
    END d4
    PIN d5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  26.30 2.62 26.72 3.26 ;
        END
    END d5
    PIN d6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  18.72 2.62 19.16 3.26 ;
        END
    END d6
    PIN d7
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  19.62 2.72 20.32 3.26 ;
        END
    END d7
    PIN sl0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.56 3.04 13.68 3.04 13.68 2.47 14.00 2.47 14.00 2.72
                 14.56 2.72 ;
        END
    END sl0
    PIN sl1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.98  LAYER metal1  ;
        ANTENNAGATEAREA 2.11  LAYER metal2  ;
        ANTENNAMAXAREACAR 0.08  LAYER metal1  ;
        ANTENNAMAXAREACAR 0.39  LAYER metal2  ;
        PORT
        LAYER metal2 ;
                POLYGON  22.36 3.90 6.76 3.90 6.76 2.74 7.08 2.74 7.08 3.58 15.76 3.58
                 15.76 2.72 16.08 2.72 16.08 3.58 22.04 3.58 22.04 2.72
                 22.36 2.72 ;
        LAYER v1 ;
        RECT  22.04 2.72 22.36 3.04 ;
        RECT  15.76 2.72 16.08 3.04 ;
        RECT  6.76 2.74 7.08 3.06 ;
        LAYER metal1 ;
        RECT  22.04 2.35 22.36 3.04 ;
        RECT  15.52 2.72 16.08 3.26 ;
        RECT  6.76 2.37 7.08 3.06 ;
        END
    END sl1
    PIN sl2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.18  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  32.02 3.68 31.52 3.68 31.52 3.36 31.70 3.36 31.70 2.62
                 32.02 2.62 ;
        END
    END sl2
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  40.80 4.32 40.46 4.32 40.46 4.00 40.48 4.00 40.48 1.66
                 40.46 1.66 40.46 1.34 40.80 1.34 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  40.96 0.90 27.00 0.90 27.00 1.14 26.68 1.14 26.68 0.90
                 19.54 0.90 19.54 1.14 19.22 1.14 19.22 0.90 16.08 0.90
                 16.08 1.14 15.76 1.14 15.76 0.90 14.00 0.90 14.00 1.14
                 13.68 1.14 13.68 0.90 10.54 0.90 10.54 1.14 10.22 1.14
                 10.22 0.90 2.98 0.90 2.98 1.14 2.66 1.14 2.66 0.90 0.00 0.90
                 0.00 -0.90 40.96 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  40.96 6.66 0.00 6.66 0.00 4.86 13.68 4.86 13.68 4.62
                 14.00 4.62 14.00 4.86 15.76 4.86 15.76 4.62 16.08 4.62
                 16.08 4.86 40.96 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  40.16 2.68 39.40 2.68 39.40 4.48 39.08 4.48 39.08 1.33
                 39.40 1.33 39.40 2.36 40.16 2.36 ;
        RECT  38.44 1.44 38.76 2.15 ;
        POLYGON  38.36 4.39 37.69 4.39 37.69 4.07 38.04 4.07 38.04 2.94
                 36.73 2.94 36.73 2.62 37.70 2.62 37.70 1.22 38.02 1.22
                 38.02 2.62 38.36 2.62 ;
        RECT  37.17 3.26 37.72 3.75 ;
        POLYGON  36.41 3.82 35.00 3.82 35.00 4.54 32.62 4.54 32.62 4.22
                 34.68 4.22 34.68 3.50 36.09 3.50 36.09 2.18 34.68 2.18
                 34.68 1.44 35.00 1.44 35.00 1.86 36.41 1.86 ;
        RECT  35.38 1.22 36.38 1.54 ;
        RECT  35.38 4.14 36.38 4.46 ;
        POLYGON  35.77 2.94 33.62 2.94 33.62 3.90 33.30 3.90 33.30 2.44
                 32.32 2.44 32.32 2.12 33.30 2.12 33.30 1.22 33.62 1.22
                 33.62 2.62 35.77 2.62 ;
        RECT  32.56 1.22 32.94 1.80 ;
        RECT  31.24 1.22 32.24 1.54 ;
        RECT  31.24 4.14 32.24 4.46 ;
        POLYGON  31.16 3.08 29.92 3.08 29.92 4.06 29.60 4.06 29.60 1.22
                 29.92 1.22 29.92 2.76 30.84 2.76 30.84 2.62 31.16 2.62 ;
        RECT  30.24 1.22 30.56 2.44 ;
        POLYGON  29.24 3.90 25.14 3.90 25.14 4.54 21.98 4.54 21.98 4.22
                 24.82 4.22 24.82 3.58 29.24 3.58 ;
        POLYGON  29.08 2.18 24.60 2.18 24.60 1.78 23.38 1.78 23.38 1.46
                 24.92 1.46 24.92 1.86 28.76 1.86 28.76 1.46 29.08 1.46 ;
        RECT  27.52 4.22 28.54 4.54 ;
        RECT  27.38 1.22 28.38 1.54 ;
        RECT  28.06 2.50 28.38 3.14 ;
        RECT  25.46 4.22 26.46 4.54 ;
        RECT  25.30 1.22 26.30 1.54 ;
        RECT  25.46 2.62 25.78 3.26 ;
        RECT  24.18 3.22 24.50 3.90 ;
        RECT  17.14 3.58 23.86 3.90 ;
        POLYGON  23.08 3.25 22.68 3.25 22.68 1.58 23.00 1.58 23.00 2.93
                 23.08 2.93 ;
        POLYGON  22.30 1.78 21.62 1.78 21.62 2.18 17.14 2.18 17.14 1.46
                 17.46 1.46 17.46 1.86 21.30 1.86 21.30 1.46 22.30 1.46 ;
        RECT  20.90 2.62 21.22 3.26 ;
        RECT  19.92 1.22 20.92 1.54 ;
        RECT  19.92 4.22 20.92 4.54 ;
        RECT  17.84 1.22 18.84 1.54 ;
        RECT  17.82 4.22 18.84 4.54 ;
        RECT  18.00 2.62 18.32 3.26 ;
        POLYGON  16.78 4.54 16.46 4.54 16.46 4.30 15.38 4.30 15.38 4.54
                 15.06 4.54 15.06 3.98 16.46 3.98 16.46 1.90 15.06 1.90
                 15.06 1.58 16.78 1.58 ;
        POLYGON  14.70 1.90 13.30 1.90 13.30 3.38 14.70 3.38 14.70 3.70
                 12.98 3.70 12.98 1.44 13.30 1.44 13.30 1.58 14.70 1.58 ;
        POLYGON  12.62 2.18 7.50 2.18 7.50 1.78 6.82 1.78 6.82 1.46 7.82 1.46
                 7.82 1.86 12.30 1.86 12.30 1.46 12.62 1.46 ;
        POLYGON  12.62 3.90 7.82 3.90 7.82 4.54 5.25 4.54 5.25 4.22 7.50 4.22
                 7.50 3.58 12.62 3.58 ;
        RECT  10.92 4.22 11.94 4.54 ;
        RECT  10.92 1.22 11.92 1.54 ;
        RECT  11.44 2.61 11.76 3.26 ;
        RECT  8.20 1.22 9.84 1.54 ;
        RECT  8.20 4.22 9.84 4.54 ;
        RECT  7.80 2.50 8.12 3.14 ;
        POLYGON  7.14 3.90 0.42 3.90 0.42 3.58 6.82 3.58 6.82 3.38 7.14 3.38 ;
        POLYGON  6.44 3.26 6.12 3.26 6.12 3.25 6.04 3.25 6.04 2.93 6.12 2.93
                 6.12 1.22 6.44 1.22 ;
        POLYGON  5.74 1.78 5.06 1.78 5.06 2.18 0.58 2.18 0.58 1.46 0.90 1.46
                 0.90 1.86 4.74 1.86 4.74 1.46 5.74 1.46 ;
        RECT  5.08 2.90 5.72 3.22 ;
        RECT  4.15 2.64 4.50 3.25 ;
        RECT  3.36 1.22 4.36 1.54 ;
        RECT  3.20 4.22 4.20 4.54 ;
        RECT  1.28 1.22 2.28 1.54 ;
        RECT  1.12 4.22 2.14 4.54 ;
        RECT  1.28 2.50 1.60 3.14 ;
        LAYER v1 ;
        RECT  38.44 1.44 38.76 1.76 ;
        RECT  37.40 3.26 37.72 3.58 ;
        RECT  34.68 1.44 35.00 1.76 ;
        RECT  32.62 1.44 32.94 1.76 ;
        RECT  30.24 1.22 30.56 1.54 ;
        RECT  28.06 2.50 28.38 2.82 ;
        RECT  25.46 2.64 25.78 2.96 ;
        RECT  24.18 3.58 24.50 3.90 ;
        RECT  22.68 2.72 23.00 3.04 ;
        RECT  20.90 2.64 21.22 2.96 ;
        RECT  18.00 2.64 18.32 2.96 ;
        RECT  16.46 4.22 16.78 4.54 ;
        RECT  15.06 4.22 15.38 4.54 ;
        RECT  12.98 1.86 13.30 2.18 ;
        RECT  11.44 2.66 11.76 2.98 ;
        RECT  7.80 2.66 8.12 2.98 ;
        RECT  6.12 1.22 6.44 1.54 ;
        RECT  5.40 2.90 5.72 3.22 ;
        RECT  4.18 2.64 4.50 2.96 ;
        RECT  1.28 2.50 1.60 2.82 ;
        LAYER metal2 ;
        RECT  32.62 1.44 38.76 1.76 ;
        POLYGON  37.72 4.32 24.82 4.32 24.82 3.04 22.68 3.04 22.68 2.72
                 25.14 2.72 25.14 4.00 37.40 4.00 37.40 3.26 37.72 3.26 ;
        RECT  6.12 1.22 30.56 1.54 ;
        POLYGON  28.38 2.82 28.06 2.82 28.06 2.18 25.78 2.18 25.78 2.96
                 25.46 2.96 25.46 2.18 21.22 2.18 21.22 2.96 20.90 2.96
                 20.90 2.18 18.32 2.18 18.32 2.96 18.00 2.96 18.00 2.18
                 11.76 2.18 11.76 2.98 11.44 2.98 11.44 2.18 8.12 2.18
                 8.12 2.98 7.80 2.98 7.80 2.18 4.50 2.18 4.50 2.96 4.18 2.96
                 4.18 2.18 1.60 2.18 1.60 2.82 1.28 2.82 1.28 1.86 28.38 1.86 ;
        POLYGON  24.50 4.54 5.40 4.54 5.40 2.90 5.72 2.90 5.72 4.22 24.18 4.22
                 24.18 3.58 24.50 3.58 ;
    END
END muxi8_1

MACRO muxi4_4
    CLASS CORE ;
    FOREIGN muxi4_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.20 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  14.05 2.08 14.56 2.62 ;
        END
    END d0
    PIN d1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  14.88 1.98 15.20 2.62 ;
        END
    END d1
    PIN d2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.15 2.60 1.76 3.04 ;
        END
    END d2
    PIN d3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.60 0.83 3.04 ;
        END
    END d3
    PIN sl0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.80  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.26 2.50 3.68 3.04 ;
        END
    END sl0
    PIN sl1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.44 3.68 8.93 3.68 8.93 2.90 9.25 2.90 9.25 3.36 9.44 3.36 ;
        END
    END sl1
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  19.04 2.40 18.80 2.40 18.80 4.54 18.48 4.54 18.48 3.98
                 17.40 3.98 17.40 4.54 17.08 4.54 17.08 3.66 18.48 3.66
                 18.48 2.14 17.08 2.14 17.08 1.22 17.40 1.22 17.40 1.82
                 18.48 1.82 18.48 1.22 18.80 1.22 18.80 2.08 19.04 2.08 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  19.20 0.90 18.10 0.90 18.10 1.50 17.78 1.50 17.78 0.90
                 16.02 0.90 16.02 1.50 15.70 1.50 15.70 0.90 1.20 0.90
                 1.20 1.54 0.88 1.54 0.88 0.90 0.00 0.90 0.00 -0.90 19.20 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  19.20 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 14.11 4.86 14.11 4.22 14.43 4.22 14.43 4.86
                 15.70 4.86 15.70 4.34 16.02 4.34 16.02 4.86 17.78 4.86
                 17.78 4.38 18.10 4.38 18.10 4.86 19.20 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  18.10 2.98 16.72 2.98 16.72 4.54 16.40 4.54 16.40 1.22
                 16.72 1.22 16.72 2.66 18.10 2.66 ;
        POLYGON  16.01 3.26 10.08 3.26 10.08 4.54 5.04 4.54 5.04 3.04 4.42 3.04
                 4.42 2.34 4.74 2.34 4.74 2.72 5.36 2.72 5.36 4.22 9.76 4.22
                 9.76 2.82 9.67 2.82 9.67 2.50 10.08 2.50 10.08 2.94 15.69 2.94
                 15.69 2.66 16.01 2.66 ;
        RECT  11.13 1.22 15.34 1.54 ;
        POLYGON  15.34 4.54 15.02 4.54 15.02 3.90 12.53 3.90 12.53 3.58
                 15.34 3.58 ;
        RECT  12.53 1.86 13.73 2.18 ;
        RECT  11.13 4.22 13.53 4.54 ;
        POLYGON  12.15 2.18 5.52 2.18 5.52 2.34 5.20 2.34 5.20 1.86 12.15 1.86 ;
        POLYGON  12.15 3.90 10.77 3.90 10.77 4.54 10.45 4.54 10.45 3.58
                 12.15 3.58 ;
        RECT  2.96 1.22 10.77 1.54 ;
        POLYGON  8.61 3.90 5.68 3.90 5.68 3.58 8.12 3.58 8.12 2.50 8.44 2.50
                 8.44 3.58 8.61 3.58 ;
        POLYGON  7.76 3.26 6.02 3.26 6.02 2.94 7.44 2.94 7.44 2.50 7.76 2.50 ;
        POLYGON  4.72 4.36 4.40 4.36 4.40 3.90 2.96 3.90 2.96 3.58 4.72 3.58 ;
        POLYGON  4.06 2.18 0.18 2.18 0.18 1.76 0.50 1.76 0.50 1.86 4.06 1.86 ;
        RECT  1.58 4.22 3.98 4.54 ;
        RECT  1.58 1.22 2.58 1.54 ;
        POLYGON  2.58 3.90 0.50 3.90 0.50 4.54 0.18 4.54 0.18 3.58 2.58 3.58 ;
    END
END muxi4_4

MACRO muxi4_2
    CLASS CORE ;
    FOREIGN muxi4_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 17.92 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  14.05 2.08 14.56 2.62 ;
        END
    END d0
    PIN d1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  14.88 1.98 15.20 2.62 ;
        END
    END d1
    PIN d2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.15 2.60 1.76 3.04 ;
        END
    END d2
    PIN d3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.60 0.83 3.04 ;
        END
    END d3
    PIN sl0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.80  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.26 2.50 3.68 3.04 ;
        END
    END sl0
    PIN sl1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.44 3.68 8.93 3.68 8.93 2.90 9.25 2.90 9.25 3.36 9.44 3.36 ;
        END
    END sl1
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  17.76 3.98 17.42 3.98 17.42 4.54 17.10 4.54 17.10 3.66
                 17.44 3.66 17.44 1.54 17.10 1.54 17.10 1.22 17.76 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  17.92 0.90 1.20 0.90 1.20 1.54 0.88 1.54 0.88 0.90 0.00 0.90
                 0.00 -0.90 17.92 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  17.92 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 14.11 4.86 14.11 4.22 14.43 4.22 14.43 4.86
                 16.40 4.86 16.40 4.34 16.72 4.34 16.72 4.86 17.92 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  16.88 3.40 16.30 3.98 16.02 3.98 16.02 4.54 15.70 4.54
                 15.70 3.66 16.16 3.66 16.56 3.26 16.56 2.22 15.88 1.54
                 15.70 1.54 15.70 1.22 16.02 1.22 16.88 2.08 ;
        POLYGON  16.08 3.26 10.08 3.26 10.08 4.54 5.04 4.54 5.04 3.04 4.42 3.04
                 4.42 2.34 4.74 2.34 4.74 2.72 5.36 2.72 5.36 4.22 9.76 4.22
                 9.76 2.82 9.67 2.82 9.67 2.50 10.08 2.50 10.08 2.94 15.76 2.94
                 15.76 2.66 16.08 2.66 ;
        RECT  11.13 1.22 15.34 1.54 ;
        POLYGON  15.34 4.54 15.02 4.54 15.02 3.90 12.53 3.90 12.53 3.58
                 15.34 3.58 ;
        RECT  12.53 1.86 13.73 2.18 ;
        RECT  11.13 4.22 13.53 4.54 ;
        POLYGON  12.15 2.18 5.52 2.18 5.52 2.34 5.20 2.34 5.20 1.86 12.15 1.86 ;
        POLYGON  12.15 3.90 10.77 3.90 10.77 4.54 10.45 4.54 10.45 3.58
                 12.15 3.58 ;
        RECT  2.96 1.22 10.77 1.54 ;
        POLYGON  8.61 3.90 5.68 3.90 5.68 3.58 8.12 3.58 8.12 2.50 8.44 2.50
                 8.44 3.58 8.61 3.58 ;
        POLYGON  7.76 3.26 6.02 3.26 6.02 2.94 7.44 2.94 7.44 2.50 7.76 2.50 ;
        POLYGON  4.72 4.36 4.40 4.36 4.40 3.90 2.96 3.90 2.96 3.58 4.72 3.58 ;
        POLYGON  4.06 2.18 0.18 2.18 0.18 1.76 0.50 1.76 0.50 1.86 4.06 1.86 ;
        RECT  1.58 4.22 3.98 4.54 ;
        RECT  1.58 1.22 2.58 1.54 ;
        POLYGON  2.58 3.90 0.50 3.90 0.50 4.54 0.18 4.54 0.18 3.58 2.58 3.58 ;
    END
END muxi4_2

MACRO muxi4_1
    CLASS CORE ;
    FOREIGN muxi4_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 17.92 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  14.05 2.08 14.56 2.62 ;
        END
    END d0
    PIN d1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  14.88 1.98 15.20 2.62 ;
        END
    END d1
    PIN d2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.15 2.60 1.76 3.04 ;
        END
    END d2
    PIN d3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.60 0.83 3.04 ;
        END
    END d3
    PIN sl0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.80  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.26 2.50 3.68 3.04 ;
        END
    END sl0
    PIN sl1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.44 3.68 8.93 3.68 8.93 2.90 9.25 2.90 9.25 3.36 9.44 3.36 ;
        END
    END sl1
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  17.76 4.54 17.10 4.54 17.10 4.22 17.44 4.22 17.44 1.54
                 17.10 1.54 17.10 1.22 17.76 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  17.92 0.90 1.20 0.90 1.20 1.54 0.88 1.54 0.88 0.90 0.00 0.90
                 0.00 -0.90 17.92 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  17.92 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 14.11 4.86 14.11 4.22 14.43 4.22 14.43 4.86
                 16.40 4.86 16.40 4.34 16.72 4.34 16.72 4.86 17.92 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  16.88 3.40 16.02 4.26 16.02 4.54 15.70 4.54 15.70 4.12
                 16.56 3.26 16.56 2.22 15.88 1.54 15.70 1.54 15.70 1.22
                 16.02 1.22 16.88 2.08 ;
        POLYGON  16.08 3.26 10.08 3.26 10.08 4.54 5.04 4.54 5.04 3.04 4.42 3.04
                 4.42 2.34 4.74 2.34 4.74 2.72 5.36 2.72 5.36 4.22 9.76 4.22
                 9.76 2.82 9.67 2.82 9.67 2.50 10.08 2.50 10.08 2.94 16.08 2.94 ;
        RECT  11.13 1.22 15.34 1.54 ;
        POLYGON  15.34 4.54 15.02 4.54 15.02 3.90 12.53 3.90 12.53 3.58
                 15.34 3.58 ;
        RECT  12.53 1.86 13.73 2.18 ;
        RECT  11.13 4.22 13.53 4.54 ;
        POLYGON  12.15 2.18 5.52 2.18 5.52 2.34 5.20 2.34 5.20 1.86 12.15 1.86 ;
        POLYGON  12.15 3.90 10.77 3.90 10.77 4.54 10.45 4.54 10.45 3.58
                 12.15 3.58 ;
        RECT  2.96 1.22 10.77 1.54 ;
        POLYGON  8.61 3.90 5.68 3.90 5.68 3.58 8.12 3.58 8.12 2.50 8.44 2.50
                 8.44 3.58 8.61 3.58 ;
        POLYGON  7.76 3.26 6.02 3.26 6.02 2.94 7.44 2.94 7.44 2.50 7.76 2.50 ;
        POLYGON  4.72 4.36 4.40 4.36 4.40 3.90 2.96 3.90 2.96 3.58 4.72 3.58 ;
        POLYGON  4.06 2.18 0.18 2.18 0.18 1.76 0.50 1.76 0.50 1.86 4.06 1.86 ;
        RECT  1.58 4.22 3.98 4.54 ;
        RECT  1.58 1.22 2.58 1.54 ;
        POLYGON  2.58 3.90 0.50 3.90 0.50 4.54 0.18 4.54 0.18 3.58 2.58 3.58 ;
    END
END muxi4_1

MACRO muxi2_4
    CLASS CORE ;
    FOREIGN muxi2_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.24 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 1.98 5.60 2.62 ;
        END
    END d0
    PIN d1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.92 1.98 6.24 2.62 ;
        END
    END d1
    PIN sl0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.17  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.40 1.12 3.04 ;
        END
    END sl0
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.08 2.40 9.95 2.40 9.95 4.54 9.63 4.54 9.63 3.90 8.55 3.90
                 8.55 4.54 8.23 4.54 8.23 3.58 9.63 3.58 9.63 2.06 8.23 2.06
                 8.23 1.22 8.55 1.22 8.55 1.74 9.63 1.74 9.63 1.22 9.95 1.22
                 9.95 2.08 10.08 2.08 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  10.24 0.90 9.25 0.90 9.25 1.42 8.93 1.42 8.93 0.90 7.17 0.90
                 7.17 1.42 6.85 1.42 6.85 0.90 1.20 0.90 1.20 1.00 0.88 1.00
                 0.88 0.90 0.00 0.90 0.00 -0.90 10.24 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  10.24 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.34 1.20 4.34
                 1.20 4.86 5.26 4.86 5.26 4.34 5.58 4.34 5.58 4.86 6.85 4.86
                 6.85 4.38 7.17 4.38 7.17 4.86 8.93 4.86 8.93 4.38 9.25 4.38
                 9.25 4.86 10.24 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  9.23 2.98 7.87 2.98 7.87 4.54 7.55 4.54 7.55 1.22 7.87 1.22
                 7.87 2.66 9.23 2.66 ;
        POLYGON  7.16 2.98 6.88 2.98 6.88 3.26 3.34 3.26 3.22 3.38 3.22 3.58
                 2.34 3.58 2.34 3.26 2.88 3.26 3.06 3.08 3.06 2.18 2.39 2.18
                 2.39 1.86 3.38 1.86 3.38 2.94 6.56 2.94 6.56 2.66 7.16 2.66 ;
        POLYGON  6.49 1.54 1.88 1.54 1.88 2.18 1.56 2.18 1.56 1.22 6.49 1.22 ;
        POLYGON  6.49 4.54 6.17 4.54 6.17 3.90 3.68 3.90 3.68 3.58 6.49 3.58 ;
        RECT  3.76 1.86 4.88 2.18 ;
        RECT  1.56 4.22 4.68 4.54 ;
        POLYGON  2.74 2.94 2.02 2.94 2.02 3.90 0.50 3.90 0.50 4.06 0.16 4.06
                 0.16 1.44 0.50 1.44 0.50 1.76 0.48 1.76 0.48 3.58 1.70 3.58
                 1.70 2.62 2.74 2.62 ;
    END
END muxi2_4

MACRO muxi2_2
    CLASS CORE ;
    FOREIGN muxi2_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.96 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 1.98 5.60 2.62 ;
        END
    END d0
    PIN d1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.92 1.98 6.24 2.62 ;
        END
    END d1
    PIN sl0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.17  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.72 1.44 3.04 ;
        END
    END sl0
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.80 3.90 8.65 3.90 8.65 4.54 8.33 4.54 8.33 3.58 8.48 3.58
                 8.48 1.54 8.33 1.54 8.33 1.22 8.80 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.96 0.90 1.20 0.90 1.20 1.00 0.88 1.00 0.88 0.90 0.00 0.90
                 0.00 -0.90 8.96 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  8.96 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.34 1.20 4.34
                 1.20 4.86 5.34 4.86 5.34 4.34 5.66 4.34 5.66 4.86 7.63 4.86
                 7.63 4.34 7.95 4.34 7.95 4.86 8.96 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  8.11 3.28 7.25 4.14 7.25 4.46 6.93 4.46 6.93 4.00 7.79 3.14
                 7.79 1.92 7.41 1.54 6.93 1.54 6.93 1.22 7.55 1.22 8.11 1.78 ;
        POLYGON  7.21 3.26 3.38 3.26 3.38 3.42 3.06 3.42 3.06 2.18 2.39 2.18
                 2.39 1.86 3.38 1.86 3.38 2.94 6.89 2.94 6.89 2.66 7.21 2.66 ;
        POLYGON  6.57 1.54 1.88 1.54 1.88 2.18 1.56 2.18 1.56 1.22 6.57 1.22 ;
        POLYGON  6.57 4.46 6.25 4.46 6.25 3.90 3.76 3.90 3.76 3.58 6.57 3.58 ;
        RECT  3.76 1.86 4.96 2.18 ;
        RECT  1.56 4.22 4.76 4.54 ;
        POLYGON  2.74 3.90 0.50 3.90 0.50 4.06 0.16 4.06 0.16 1.44 0.50 1.44
                 0.50 1.76 0.48 1.76 0.48 3.58 2.42 3.58 2.42 2.62 2.74 2.62 ;
    END
END muxi2_2

MACRO muxi2_1
    CLASS CORE ;
    FOREIGN muxi2_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.96 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 1.98 5.60 2.62 ;
        END
    END d0
    PIN d1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.92 1.98 6.24 2.62 ;
        END
    END d1
    PIN sl0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.17  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.72 1.44 3.04 ;
        END
    END sl0
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.80 4.06 8.33 4.06 8.33 3.74 8.48 3.74 8.48 1.54 8.33 1.54
                 8.33 1.22 8.80 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.96 0.90 1.20 0.90 1.20 1.00 0.88 1.00 0.88 0.90 0.00 0.90
                 0.00 -0.90 8.96 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  8.96 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.34 1.20 4.34
                 1.20 4.86 5.34 4.86 5.34 4.34 5.66 4.34 5.66 4.86 7.63 4.86
                 7.63 4.34 7.95 4.34 7.95 4.86 8.96 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  8.11 3.28 7.25 4.14 7.25 4.46 6.93 4.46 6.93 4.00 7.79 3.14
                 7.79 1.92 7.41 1.54 6.93 1.54 6.93 1.22 7.55 1.22 8.11 1.78 ;
        POLYGON  7.21 3.26 3.38 3.26 3.38 3.42 3.06 3.42 3.06 2.18 2.39 2.18
                 2.39 1.86 3.38 1.86 3.38 2.94 7.21 2.94 ;
        POLYGON  6.57 1.54 1.88 1.54 1.88 2.18 1.56 2.18 1.56 1.22 6.57 1.22 ;
        POLYGON  6.57 4.46 6.25 4.46 6.25 3.90 3.76 3.90 3.76 3.58 6.57 3.58 ;
        RECT  3.76 1.86 4.96 2.18 ;
        RECT  1.56 4.22 4.76 4.54 ;
        POLYGON  2.74 3.90 0.50 3.90 0.50 4.06 0.16 4.06 0.16 1.44 0.50 1.44
                 0.50 1.76 0.48 1.76 0.48 3.58 2.42 3.58 2.42 2.62 2.74 2.62 ;
    END
END muxi2_1

MACRO mux8_4
    CLASS CORE ;
    FOREIGN mux8_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 40.32 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.62 2.52 3.26 ;
        END
    END d0
    PIN d1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.96 2.72 3.68 3.12 ;
        END
    END d1
    PIN d2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.40 2.72 10.94 3.16 ;
        END
    END d2
    PIN d3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  9.12 2.54 9.44 3.18 ;
        END
    END d3
    PIN d4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  27.04 2.63 27.50 3.26 ;
        END
    END d4
    PIN d5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  26.34 2.62 26.72 3.26 ;
        END
    END d5
    PIN d6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  18.72 2.62 19.16 3.26 ;
        END
    END d6
    PIN d7
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  19.62 2.72 20.32 3.26 ;
        END
    END d7
    PIN sl0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.56 3.04 13.68 3.04 13.68 2.47 14.00 2.47 14.00 2.72
                 14.56 2.72 ;
        END
    END sl0
    PIN sl1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.98  LAYER metal1  ;
        ANTENNAGATEAREA 2.11  LAYER metal2  ;
        ANTENNAMAXAREACAR 0.02  LAYER metal1  ;
        ANTENNAMAXAREACAR 0.39  LAYER metal2  ;
        PORT
        LAYER metal2 ;
                POLYGON  22.36 3.90 6.76 3.90 6.76 2.74 7.08 2.74 7.08 3.58 15.76 3.58
                 15.76 2.72 16.08 2.72 16.08 3.58 22.04 3.58 22.04 2.72
                 22.36 2.72 ;
        LAYER v1 ;
        RECT  22.04 2.72 22.36 3.04 ;
        RECT  15.76 2.72 16.08 3.04 ;
        RECT  6.76 2.74 7.08 3.06 ;
        LAYER metal1 ;
        RECT  22.04 2.35 22.36 3.04 ;
        RECT  15.52 2.62 16.08 3.26 ;
        RECT  6.76 2.37 7.08 3.06 ;
        END
    END sl1
    PIN sl2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.18  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  32.06 3.68 31.52 3.68 31.52 3.36 31.74 3.36 31.74 2.62
                 32.06 2.62 ;
        END
    END sl2
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  40.16 4.54 38.42 4.54 38.42 4.22 39.84 4.22 39.84 1.54
                 38.42 1.54 38.42 1.22 40.16 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  40.32 0.90 27.04 0.90 27.04 1.14 26.72 1.14 26.72 0.90
                 19.54 0.90 19.54 1.14 19.22 1.14 19.22 0.90 16.08 0.90
                 16.08 1.14 15.76 1.14 15.76 0.90 14.00 0.90 14.00 1.14
                 13.68 1.14 13.68 0.90 10.54 0.90 10.54 1.14 10.22 1.14
                 10.22 0.90 2.98 0.90 2.98 1.14 2.66 1.14 2.66 0.90 0.00 0.90
                 0.00 -0.90 40.32 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  40.32 6.66 0.00 6.66 0.00 4.86 13.68 4.86 13.68 4.62
                 14.00 4.62 14.00 4.86 15.76 4.86 15.76 4.62 16.08 4.62
                 16.08 4.86 40.32 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  39.12 1.91 39.44 2.74 ;
        POLYGON  38.42 3.90 37.73 3.90 37.73 3.58 38.10 3.58 38.10 2.62
                 36.52 2.62 36.52 2.30 37.74 2.30 37.74 1.22 38.06 1.22
                 38.06 2.30 38.42 2.30 ;
        RECT  37.15 2.94 37.78 3.26 ;
        RECT  35.42 1.22 36.42 1.54 ;
        RECT  35.42 4.14 36.42 4.46 ;
        POLYGON  35.21 3.82 35.04 3.82 35.04 4.54 32.66 4.54 32.66 4.22
                 34.72 4.22 34.72 3.50 34.89 3.50 34.89 2.18 34.72 2.18
                 34.72 1.44 35.04 1.44 35.04 1.86 35.21 1.86 ;
        POLYGON  34.57 3.04 33.66 3.04 33.66 3.90 33.34 3.90 33.34 2.44
                 32.36 2.44 32.36 2.12 33.34 2.12 33.34 1.22 33.66 1.22
                 33.66 2.72 34.57 2.72 ;
        RECT  32.60 1.22 32.98 1.80 ;
        RECT  31.28 1.22 32.28 1.54 ;
        RECT  31.28 4.14 32.28 4.46 ;
        POLYGON  31.20 3.08 29.96 3.08 29.96 4.06 29.64 4.06 29.64 1.22
                 29.96 1.22 29.96 2.76 30.88 2.76 30.88 2.62 31.20 2.62 ;
        RECT  30.28 1.22 30.60 2.44 ;
        POLYGON  29.28 3.90 25.14 3.90 25.14 4.54 21.98 4.54 21.98 4.22
                 24.82 4.22 24.82 3.58 29.28 3.58 ;
        POLYGON  29.12 2.18 24.64 2.18 24.64 1.78 23.38 1.78 23.38 1.46
                 24.96 1.46 24.96 1.86 28.80 1.86 28.80 1.46 29.12 1.46 ;
        RECT  27.56 4.22 28.58 4.54 ;
        RECT  27.42 1.22 28.42 1.54 ;
        RECT  28.10 2.50 28.42 3.14 ;
        RECT  25.50 4.22 26.50 4.54 ;
        RECT  25.34 1.22 26.34 1.54 ;
        RECT  25.46 2.52 25.78 3.26 ;
        RECT  24.18 3.04 24.50 3.68 ;
        RECT  17.14 3.58 23.86 3.90 ;
        POLYGON  23.08 3.25 22.68 3.25 22.68 1.58 23.00 1.58 23.00 2.93
                 23.08 2.93 ;
        POLYGON  22.30 1.78 21.62 1.78 21.62 2.18 17.14 2.18 17.14 1.46
                 17.46 1.46 17.46 1.86 21.30 1.86 21.30 1.46 22.30 1.46 ;
        RECT  20.90 2.62 21.22 3.26 ;
        RECT  19.92 1.22 20.92 1.54 ;
        RECT  19.92 4.22 20.92 4.54 ;
        RECT  17.84 1.22 18.84 1.54 ;
        RECT  17.82 4.22 18.84 4.54 ;
        RECT  18.00 2.62 18.32 3.26 ;
        POLYGON  16.79 4.54 16.47 4.54 16.47 4.30 15.38 4.30 15.38 4.54
                 15.06 4.54 15.06 3.98 16.47 3.98 16.47 1.90 15.06 1.90
                 15.06 1.58 16.79 1.58 ;
        POLYGON  14.70 1.90 13.30 1.90 13.30 3.38 14.70 3.38 14.70 3.70
                 12.98 3.70 12.98 1.44 13.30 1.44 13.30 1.58 14.70 1.58 ;
        POLYGON  12.62 2.18 7.50 2.18 7.50 1.78 6.82 1.78 6.82 1.46 7.82 1.46
                 7.82 1.86 12.30 1.86 12.30 1.46 12.62 1.46 ;
        POLYGON  12.62 3.90 7.82 3.90 7.82 4.54 5.25 4.54 5.25 4.22 7.50 4.22
                 7.50 3.58 12.62 3.58 ;
        RECT  10.92 4.22 11.94 4.54 ;
        RECT  10.92 1.22 11.92 1.54 ;
        RECT  11.44 2.61 11.76 3.26 ;
        RECT  8.20 1.22 9.84 1.54 ;
        RECT  8.20 4.22 9.84 4.54 ;
        RECT  7.80 2.50 8.12 3.14 ;
        POLYGON  7.14 3.90 0.42 3.90 0.42 3.58 6.82 3.58 6.82 3.38 7.14 3.38 ;
        POLYGON  6.44 3.26 6.12 3.26 6.12 3.25 6.04 3.25 6.04 2.93 6.12 2.93
                 6.12 1.22 6.44 1.22 ;
        POLYGON  5.74 1.78 5.06 1.78 5.06 2.18 0.58 2.18 0.58 1.46 0.90 1.46
                 0.90 1.86 4.74 1.86 4.74 1.46 5.74 1.46 ;
        RECT  5.08 2.90 5.72 3.22 ;
        RECT  4.15 2.64 4.50 3.25 ;
        RECT  3.36 1.22 4.36 1.54 ;
        RECT  3.20 4.22 4.20 4.54 ;
        RECT  1.28 1.22 2.28 1.54 ;
        RECT  1.12 4.22 2.14 4.54 ;
        RECT  1.28 2.50 1.60 3.14 ;
        LAYER v1 ;
        RECT  39.12 1.91 39.44 2.23 ;
        RECT  37.46 2.94 37.78 3.26 ;
        RECT  34.72 1.44 35.04 1.76 ;
        RECT  32.66 1.44 32.98 1.76 ;
        RECT  30.28 1.22 30.60 1.54 ;
        RECT  28.10 2.50 28.42 2.82 ;
        RECT  25.46 2.64 25.78 2.96 ;
        RECT  24.18 3.36 24.50 3.68 ;
        RECT  22.68 2.72 23.00 3.04 ;
        RECT  20.90 2.64 21.22 2.96 ;
        RECT  18.00 2.64 18.32 2.96 ;
        RECT  16.47 4.22 16.79 4.54 ;
        RECT  15.06 4.22 15.38 4.54 ;
        RECT  12.98 1.86 13.30 2.18 ;
        RECT  11.44 2.66 11.76 2.98 ;
        RECT  7.80 2.66 8.12 2.98 ;
        RECT  6.12 1.22 6.44 1.54 ;
        RECT  5.40 2.90 5.72 3.22 ;
        RECT  4.18 2.64 4.50 2.96 ;
        RECT  1.28 2.50 1.60 2.82 ;
        LAYER metal2 ;
        POLYGON  39.44 2.23 39.12 2.23 39.12 1.76 32.66 1.76 32.66 1.44
                 39.44 1.44 ;
        POLYGON  37.78 4.32 24.82 4.32 24.82 3.04 22.68 3.04 22.68 2.72
                 25.14 2.72 25.14 4.00 37.46 4.00 37.46 2.94 37.78 2.94 ;
        RECT  6.12 1.22 30.60 1.54 ;
        POLYGON  28.42 2.82 28.10 2.82 28.10 2.18 25.78 2.18 25.78 2.96
                 25.46 2.96 25.46 2.18 21.22 2.18 21.22 2.96 20.90 2.96
                 20.90 2.18 18.32 2.18 18.32 2.96 18.00 2.96 18.00 2.18
                 11.76 2.18 11.76 2.98 11.44 2.98 11.44 2.18 8.12 2.18
                 8.12 2.98 7.80 2.98 7.80 2.18 4.50 2.18 4.50 2.96 4.18 2.96
                 4.18 2.18 1.60 2.18 1.60 2.82 1.28 2.82 1.28 1.86 28.42 1.86 ;
        POLYGON  24.50 4.54 5.40 4.54 5.40 2.90 5.72 2.90 5.72 4.22 24.18 4.22
                 24.18 3.36 24.50 3.36 ;
    END
END mux8_4

MACRO mux8_2
    CLASS CORE ;
    FOREIGN mux8_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 39.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.62 2.52 3.26 ;
        END
    END d0
    PIN d1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.96 2.72 3.68 3.12 ;
        END
    END d1
    PIN d2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.40 2.72 10.94 3.16 ;
        END
    END d2
    PIN d3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  9.12 2.54 9.44 3.18 ;
        END
    END d3
    PIN d4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  27.04 2.72 27.52 3.26 ;
        END
    END d4
    PIN d5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  26.30 2.72 26.72 3.26 ;
        END
    END d5
    PIN d6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  18.72 2.62 19.16 3.26 ;
        END
    END d6
    PIN d7
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  19.62 2.72 20.32 3.26 ;
        END
    END d7
    PIN sl0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.56 3.04 13.68 3.04 13.68 2.47 14.00 2.47 14.00 2.72
                 14.56 2.72 ;
        END
    END sl0
    PIN sl1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.98  LAYER metal1  ;
        ANTENNAGATEAREA 2.11  LAYER metal2  ;
        ANTENNAMAXAREACAR 0.02  LAYER metal1  ;
        ANTENNAMAXAREACAR 0.39  LAYER metal2  ;
        PORT
        LAYER metal2 ;
                POLYGON  22.36 3.90 6.76 3.90 6.76 2.74 7.08 2.74 7.08 3.58 15.76 3.58
                 15.76 2.72 16.08 2.72 16.08 3.58 22.04 3.58 22.04 2.72
                 22.36 2.72 ;
        LAYER v1 ;
        RECT  22.04 2.72 22.36 3.04 ;
        RECT  15.76 2.72 16.08 3.04 ;
        RECT  6.76 2.74 7.08 3.06 ;
        LAYER metal1 ;
        RECT  22.04 2.35 22.36 3.04 ;
        RECT  15.52 2.62 16.08 3.26 ;
        RECT  6.76 2.37 7.08 3.06 ;
        END
    END sl1
    PIN sl2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.18  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  32.08 3.68 31.52 3.68 31.52 3.36 31.76 3.36 31.76 2.62
                 32.08 2.62 ;
        END
    END sl2
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  39.52 3.76 39.18 3.76 39.18 3.44 39.20 3.44 39.20 1.59
                 39.18 1.59 39.18 1.27 39.52 1.27 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  39.68 0.90 27.06 0.90 27.06 1.14 26.74 1.14 26.74 0.90
                 19.54 0.90 19.54 1.14 19.22 1.14 19.22 0.90 16.08 0.90
                 16.08 1.14 15.76 1.14 15.76 0.90 14.00 0.90 14.00 1.14
                 13.68 1.14 13.68 0.90 10.54 0.90 10.54 1.14 10.22 1.14
                 10.22 0.90 2.98 0.90 2.98 1.14 2.66 1.14 2.66 0.90 0.00 0.90
                 0.00 -0.90 39.68 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  39.68 6.66 0.00 6.66 0.00 4.86 13.68 4.86 13.68 4.62
                 14.00 4.62 14.00 4.86 15.76 4.86 15.76 4.62 16.08 4.62
                 16.08 4.86 39.68 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  38.56 1.76 38.88 2.45 ;
        POLYGON  38.24 4.39 37.75 4.39 37.75 4.07 37.92 4.07 37.92 3.15
                 36.64 3.15 36.64 2.62 36.96 2.62 36.96 2.83 37.92 2.83
                 37.92 1.54 37.76 1.54 37.76 1.22 38.24 1.22 ;
        RECT  37.24 1.86 37.60 2.44 ;
        RECT  35.44 1.22 36.44 1.54 ;
        RECT  35.44 4.14 36.44 4.46 ;
        POLYGON  35.22 3.82 35.06 3.82 35.06 4.54 32.68 4.54 32.68 4.22
                 34.74 4.22 34.74 3.50 34.90 3.50 34.90 2.18 34.74 2.18
                 34.74 1.44 35.06 1.44 35.06 1.86 35.22 1.86 ;
        POLYGON  34.58 3.04 33.68 3.04 33.68 3.90 33.36 3.90 33.36 2.44
                 32.38 2.44 32.38 2.12 33.36 2.12 33.36 1.22 33.68 1.22
                 33.68 2.72 34.58 2.72 ;
        RECT  32.62 1.22 33.00 1.80 ;
        RECT  31.30 1.22 32.30 1.54 ;
        RECT  31.30 4.14 32.30 4.46 ;
        POLYGON  31.22 3.08 29.98 3.08 29.98 4.06 29.66 4.06 29.66 1.22
                 29.98 1.22 29.98 2.76 30.90 2.76 30.90 2.62 31.22 2.62 ;
        RECT  30.30 1.22 30.62 2.44 ;
        POLYGON  29.30 3.90 25.14 3.90 25.14 4.54 21.98 4.54 21.98 4.22
                 24.82 4.22 24.82 3.58 29.30 3.58 ;
        POLYGON  29.14 2.18 24.66 2.18 24.66 1.78 23.38 1.78 23.38 1.46
                 24.98 1.46 24.98 1.86 28.82 1.86 28.82 1.46 29.14 1.46 ;
        RECT  27.58 4.22 28.60 4.54 ;
        RECT  27.44 1.22 28.44 1.54 ;
        RECT  28.12 2.50 28.44 3.14 ;
        RECT  25.52 4.22 26.52 4.54 ;
        RECT  25.36 1.22 26.36 1.54 ;
        RECT  25.46 2.62 25.78 3.26 ;
        RECT  24.18 3.12 24.50 3.90 ;
        RECT  17.14 3.58 23.86 3.90 ;
        POLYGON  23.08 3.26 22.68 3.26 22.68 1.58 23.00 1.58 23.00 2.94
                 23.08 2.94 ;
        POLYGON  22.30 1.78 21.62 1.78 21.62 2.18 17.14 2.18 17.14 1.46
                 17.46 1.46 17.46 1.86 21.30 1.86 21.30 1.46 22.30 1.46 ;
        RECT  20.90 2.62 21.22 3.26 ;
        RECT  19.92 1.22 20.92 1.54 ;
        RECT  19.92 4.22 20.92 4.54 ;
        RECT  17.84 1.22 18.84 1.54 ;
        RECT  17.82 4.22 18.84 4.54 ;
        RECT  18.00 2.62 18.32 3.26 ;
        POLYGON  16.79 4.54 16.47 4.54 16.47 4.30 15.38 4.30 15.38 4.54
                 15.06 4.54 15.06 3.98 16.47 3.98 16.47 1.90 15.06 1.90
                 15.06 1.58 16.79 1.58 ;
        POLYGON  14.70 1.90 13.30 1.90 13.30 3.38 14.70 3.38 14.70 3.70
                 12.98 3.70 12.98 1.44 13.30 1.44 13.30 1.58 14.70 1.58 ;
        POLYGON  12.62 2.18 7.50 2.18 7.50 1.78 6.82 1.78 6.82 1.46 7.82 1.46
                 7.82 1.86 12.30 1.86 12.30 1.46 12.62 1.46 ;
        POLYGON  12.62 3.90 7.82 3.90 7.82 4.54 5.25 4.54 5.25 4.22 7.50 4.22
                 7.50 3.58 12.62 3.58 ;
        RECT  10.92 4.22 11.94 4.54 ;
        RECT  10.92 1.22 11.92 1.54 ;
        RECT  11.44 2.61 11.76 3.26 ;
        RECT  8.20 1.22 9.84 1.54 ;
        RECT  8.20 4.22 9.84 4.54 ;
        RECT  7.80 2.50 8.12 3.14 ;
        POLYGON  7.14 3.90 0.42 3.90 0.42 3.58 6.82 3.58 6.82 3.38 7.14 3.38 ;
        POLYGON  6.44 3.26 6.12 3.26 6.12 3.25 6.04 3.25 6.04 2.93 6.12 2.93
                 6.12 1.22 6.44 1.22 ;
        POLYGON  5.74 1.78 5.06 1.78 5.06 2.18 0.58 2.18 0.58 1.46 0.90 1.46
                 0.90 1.86 4.74 1.86 4.74 1.46 5.74 1.46 ;
        RECT  5.08 2.90 5.72 3.22 ;
        RECT  4.15 2.64 4.50 3.25 ;
        RECT  3.36 1.22 4.36 1.54 ;
        RECT  3.20 4.22 4.20 4.54 ;
        RECT  1.28 1.22 2.28 1.54 ;
        RECT  1.12 4.22 2.14 4.54 ;
        RECT  1.28 2.50 1.60 3.14 ;
        LAYER v1 ;
        RECT  38.56 1.76 38.88 2.08 ;
        RECT  37.28 2.12 37.60 2.44 ;
        RECT  34.74 1.44 35.06 1.76 ;
        RECT  32.68 1.44 33.00 1.76 ;
        RECT  30.30 1.22 30.62 1.54 ;
        RECT  28.12 2.50 28.44 2.82 ;
        RECT  25.46 2.64 25.78 2.96 ;
        RECT  24.18 3.58 24.50 3.90 ;
        RECT  22.76 2.94 23.08 3.26 ;
        RECT  20.90 2.64 21.22 2.96 ;
        RECT  18.00 2.64 18.32 2.96 ;
        RECT  16.47 4.22 16.79 4.54 ;
        RECT  15.06 4.22 15.38 4.54 ;
        RECT  12.98 1.86 13.30 2.18 ;
        RECT  11.44 2.66 11.76 2.98 ;
        RECT  7.80 2.66 8.12 2.98 ;
        RECT  6.12 1.22 6.44 1.54 ;
        RECT  5.40 2.90 5.72 3.22 ;
        RECT  4.18 2.64 4.50 2.96 ;
        RECT  1.28 2.50 1.60 2.82 ;
        LAYER metal2 ;
        POLYGON  38.88 2.08 38.56 2.08 38.56 1.76 32.68 1.76 32.68 1.44
                 38.88 1.44 ;
        POLYGON  37.60 4.32 24.82 4.32 24.82 3.26 22.76 3.26 22.76 2.94
                 25.14 2.94 25.14 4.00 37.28 4.00 37.28 2.12 37.60 2.12 ;
        RECT  6.12 1.22 30.62 1.54 ;
        POLYGON  28.44 2.82 28.12 2.82 28.12 2.18 25.78 2.18 25.78 2.96
                 25.46 2.96 25.46 2.18 21.22 2.18 21.22 2.96 20.90 2.96
                 20.90 2.18 18.32 2.18 18.32 2.96 18.00 2.96 18.00 2.18
                 11.76 2.18 11.76 2.98 11.44 2.98 11.44 2.18 8.12 2.18
                 8.12 2.98 7.80 2.98 7.80 2.18 4.50 2.18 4.50 2.96 4.18 2.96
                 4.18 2.18 1.60 2.18 1.60 2.82 1.28 2.82 1.28 1.86 28.44 1.86 ;
        POLYGON  24.50 4.54 5.40 4.54 5.40 2.90 5.72 2.90 5.72 4.22 24.18 4.22
                 24.18 3.58 24.50 3.58 ;
    END
END mux8_2

MACRO mux8_1
    CLASS CORE ;
    FOREIGN mux8_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 39.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.62 2.52 3.26 ;
        END
    END d0
    PIN d1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.96 2.72 3.68 3.12 ;
        END
    END d1
    PIN d2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.40 2.72 10.94 3.16 ;
        END
    END d2
    PIN d3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  9.12 2.54 9.44 3.18 ;
        END
    END d3
    PIN d4
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  27.18 2.72 27.66 3.15 ;
        END
    END d4
    PIN d5
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  26.30 2.72 26.86 3.15 ;
        END
    END d5
    PIN d6
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  18.72 2.62 19.14 3.26 ;
        END
    END d6
    PIN d7
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  19.62 2.72 20.32 3.06 ;
        END
    END d7
    PIN sl0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  13.68 2.72 14.56 3.04 ;
        END
    END sl0
    PIN sl1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.98  LAYER metal1  ;
        ANTENNAGATEAREA 2.11  LAYER metal2  ;
        ANTENNAMAXAREACAR 0.02  LAYER metal1  ;
        ANTENNAMAXAREACAR 0.39  LAYER metal2  ;
        PORT
        LAYER metal2 ;
                POLYGON  22.36 3.90 6.76 3.90 6.76 2.74 7.08 2.74 7.08 3.58 15.76 3.58
                 15.76 2.72 16.08 2.72 16.08 3.58 22.04 3.58 22.04 2.72
                 22.36 2.72 ;
        LAYER v1 ;
        RECT  22.04 2.72 22.36 3.04 ;
        RECT  15.76 2.72 16.08 3.04 ;
        RECT  6.76 2.74 7.08 3.06 ;
        LAYER metal1 ;
        RECT  22.04 2.35 22.36 3.04 ;
        RECT  15.52 2.62 16.08 3.26 ;
        RECT  6.76 2.37 7.08 3.06 ;
        END
    END sl1
    PIN sl2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.18  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  32.02 3.68 31.66 3.68 31.66 3.36 31.70 3.36 31.70 2.62
                 32.02 2.62 ;
        END
    END sl2
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  39.52 4.32 39.18 4.32 39.18 4.00 39.20 4.00 39.20 1.54
                 39.18 1.54 39.18 1.22 39.52 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  39.68 0.90 27.00 0.90 27.00 1.14 26.68 1.14 26.68 0.90
                 19.54 0.90 19.54 1.14 19.22 1.14 19.22 0.90 16.08 0.90
                 16.08 1.14 15.76 1.14 15.76 0.90 14.00 0.90 14.00 1.14
                 13.68 1.14 13.68 0.90 10.54 0.90 10.54 1.14 10.22 1.14
                 10.22 0.90 2.98 0.90 2.98 1.14 2.66 1.14 2.66 0.90 0.00 0.90
                 0.00 -0.90 39.68 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  39.68 6.66 0.00 6.66 0.00 4.86 13.68 4.86 13.68 4.62
                 14.00 4.62 14.00 4.86 15.76 4.86 15.76 4.62 16.08 4.62
                 16.08 4.86 39.68 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  38.54 1.44 38.86 2.07 ;
        POLYGON  38.36 4.39 37.69 4.39 37.69 4.07 38.04 4.07 38.04 2.68
                 36.73 2.68 36.73 2.36 37.70 2.36 37.70 1.22 38.02 1.22
                 38.02 2.36 38.36 2.36 ;
        RECT  37.40 3.07 37.72 3.71 ;
        POLYGON  36.41 3.82 35.00 3.82 35.00 4.54 32.62 4.54 32.62 4.22
                 34.68 4.22 34.68 3.50 36.09 3.50 36.09 2.18 34.68 2.18
                 34.68 1.44 35.00 1.44 35.00 1.86 36.41 1.86 ;
        RECT  35.38 1.22 36.38 1.54 ;
        RECT  35.38 4.14 36.38 4.46 ;
        POLYGON  35.77 2.94 33.62 2.94 33.62 3.90 33.30 3.90 33.30 2.44
                 32.32 2.44 32.32 2.12 33.30 2.12 33.30 1.22 33.62 1.22
                 33.62 2.62 35.77 2.62 ;
        RECT  32.56 1.22 32.94 1.80 ;
        RECT  31.24 1.22 32.24 1.54 ;
        RECT  31.24 4.14 32.24 4.46 ;
        POLYGON  31.16 3.08 29.92 3.08 29.92 4.06 29.60 4.06 29.60 1.22
                 29.92 1.22 29.92 2.76 30.84 2.76 30.84 2.62 31.16 2.62 ;
        RECT  30.24 1.22 30.56 2.44 ;
        POLYGON  29.24 3.90 25.14 3.90 25.14 4.54 21.98 4.54 21.98 4.22
                 24.82 4.22 24.82 3.58 29.24 3.58 ;
        POLYGON  29.08 2.18 24.60 2.18 24.60 1.54 23.38 1.54 23.38 1.22
                 24.92 1.22 24.92 1.86 28.76 1.86 28.76 1.46 29.08 1.46 ;
        RECT  27.52 4.22 28.54 4.54 ;
        RECT  27.38 1.22 28.38 1.54 ;
        RECT  28.06 2.50 28.38 3.14 ;
        RECT  25.46 4.22 26.46 4.54 ;
        RECT  25.30 1.22 26.30 1.54 ;
        RECT  25.37 2.64 25.78 3.26 ;
        RECT  24.18 3.20 24.50 3.90 ;
        RECT  17.14 3.58 23.86 3.90 ;
        POLYGON  23.08 3.26 22.68 3.26 22.68 2.00 23.00 2.00 23.00 2.94
                 23.08 2.94 ;
        POLYGON  22.30 2.00 21.62 2.00 21.62 2.18 17.14 2.18 17.14 1.46
                 17.46 1.46 17.46 1.86 21.29 1.86 21.29 1.68 22.30 1.68 ;
        RECT  20.90 2.62 21.22 3.26 ;
        RECT  19.92 1.22 20.92 1.54 ;
        RECT  19.92 4.22 20.92 4.54 ;
        RECT  17.84 1.22 18.84 1.54 ;
        RECT  17.82 4.22 18.84 4.54 ;
        RECT  18.00 2.62 18.32 3.26 ;
        POLYGON  16.78 4.54 16.46 4.54 16.46 4.30 15.38 4.30 15.38 4.54
                 15.06 4.54 15.06 3.98 16.46 3.98 16.46 1.90 15.06 1.90
                 15.06 1.58 16.78 1.58 ;
        POLYGON  14.70 1.90 13.30 1.90 13.30 3.38 14.70 3.38 14.70 3.70
                 12.98 3.70 12.98 1.58 14.70 1.58 ;
        POLYGON  12.62 2.18 7.50 2.18 7.50 1.78 6.82 1.78 6.82 1.46 7.82 1.46
                 7.82 1.86 12.30 1.86 12.30 1.46 12.62 1.46 ;
        POLYGON  12.62 3.90 7.82 3.90 7.82 4.54 5.25 4.54 5.25 4.22 7.50 4.22
                 7.50 3.58 12.62 3.58 ;
        RECT  10.92 4.22 11.94 4.54 ;
        RECT  10.92 1.22 11.92 1.54 ;
        RECT  11.44 2.61 11.76 3.26 ;
        RECT  8.20 1.22 9.84 1.54 ;
        RECT  8.20 4.22 9.84 4.54 ;
        RECT  7.80 2.50 8.12 3.14 ;
        POLYGON  7.14 3.90 0.42 3.90 0.42 3.58 6.82 3.58 6.82 3.38 7.14 3.38 ;
        POLYGON  6.44 3.26 6.12 3.26 6.12 3.25 6.04 3.25 6.04 2.93 6.12 2.93
                 6.12 1.22 6.44 1.22 ;
        POLYGON  5.74 1.78 5.06 1.78 5.06 2.18 0.58 2.18 0.58 1.46 0.90 1.46
                 0.90 1.86 4.74 1.86 4.74 1.46 5.74 1.46 ;
        RECT  5.08 2.90 5.72 3.22 ;
        RECT  4.15 2.64 4.50 3.25 ;
        RECT  3.36 1.22 4.36 1.54 ;
        RECT  3.20 4.22 4.20 4.54 ;
        RECT  1.28 1.22 2.28 1.54 ;
        RECT  1.12 4.22 2.14 4.54 ;
        RECT  1.28 2.50 1.60 3.14 ;
        LAYER v1 ;
        RECT  38.54 1.44 38.86 1.76 ;
        RECT  37.40 3.07 37.72 3.39 ;
        RECT  34.68 1.44 35.00 1.76 ;
        RECT  32.62 1.44 32.94 1.76 ;
        RECT  30.24 1.22 30.56 1.54 ;
        RECT  28.06 2.50 28.38 2.82 ;
        RECT  25.46 2.64 25.78 2.96 ;
        RECT  24.18 3.36 24.50 3.68 ;
        RECT  22.68 2.72 23.00 3.04 ;
        RECT  20.90 2.64 21.22 2.96 ;
        RECT  18.00 2.64 18.32 2.96 ;
        RECT  16.46 4.22 16.78 4.54 ;
        RECT  15.06 4.22 15.38 4.54 ;
        RECT  12.98 1.86 13.30 2.18 ;
        RECT  11.44 2.66 11.76 2.98 ;
        RECT  7.80 2.66 8.12 2.98 ;
        RECT  6.12 1.22 6.44 1.54 ;
        RECT  5.40 2.90 5.72 3.22 ;
        RECT  4.18 2.64 4.50 2.96 ;
        RECT  1.28 2.50 1.60 2.82 ;
        LAYER metal2 ;
        RECT  32.62 1.44 38.86 1.76 ;
        POLYGON  37.72 4.32 24.82 4.32 24.82 3.04 22.68 3.04 22.68 2.72
                 25.14 2.72 25.14 4.00 37.40 4.00 37.40 3.07 37.72 3.07 ;
        RECT  6.12 1.22 30.56 1.54 ;
        POLYGON  28.38 2.82 28.06 2.82 28.06 2.18 25.78 2.18 25.78 2.96
                 25.46 2.96 25.46 2.18 21.22 2.18 21.22 2.96 20.90 2.96
                 20.90 2.18 18.32 2.18 18.32 2.96 18.00 2.96 18.00 2.18
                 11.76 2.18 11.76 2.98 11.44 2.98 11.44 2.18 8.12 2.18
                 8.12 2.98 7.80 2.98 7.80 2.18 4.50 2.18 4.50 2.96 4.18 2.96
                 4.18 2.18 1.60 2.18 1.60 2.82 1.28 2.82 1.28 1.86 28.38 1.86 ;
        POLYGON  24.50 4.54 5.40 4.54 5.40 2.90 5.72 2.90 5.72 4.22 24.18 4.22
                 24.18 3.36 24.50 3.36 ;
    END
END mux8_1

MACRO mux4_4
    CLASS CORE ;
    FOREIGN mux4_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 17.92 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  14.05 2.08 14.56 2.62 ;
        END
    END d0
    PIN d1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  14.88 1.98 15.20 2.62 ;
        END
    END d1
    PIN d2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.15 2.60 1.76 3.04 ;
        END
    END d2
    PIN d3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.60 0.83 3.04 ;
        END
    END d3
    PIN sl0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.80  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.26 2.50 3.68 3.04 ;
        END
    END sl0
    PIN sl1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.44 3.68 8.93 3.68 8.93 2.90 9.25 2.90 9.25 3.36 9.44 3.36 ;
        END
    END sl1
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  17.42 4.54 17.10 4.54 17.10 3.98 16.02 3.98 16.02 4.54
                 15.70 4.54 15.70 3.66 17.10 3.66 17.10 2.40 16.80 2.40
                 16.80 2.08 17.10 2.08 17.10 1.54 15.70 1.54 15.70 1.22
                 17.42 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 17.92 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  17.92 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 14.11 4.86 14.11 4.22 14.43 4.22 14.43 4.86
                 16.40 4.86 16.40 4.30 16.72 4.30 16.72 4.86 17.92 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  16.08 3.26 10.08 3.26 10.08 4.54 5.04 4.54 5.04 3.04 4.42 3.04
                 4.42 2.34 4.74 2.34 4.74 2.72 5.36 2.72 5.36 4.22 9.76 4.22
                 9.76 2.82 9.67 2.82 9.67 2.50 10.08 2.50 10.08 2.94 15.76 2.94
                 15.76 2.62 16.08 2.62 ;
        RECT  11.13 1.22 15.34 1.54 ;
        POLYGON  15.34 4.54 15.02 4.54 15.02 3.90 12.53 3.90 12.53 3.58
                 15.34 3.58 ;
        RECT  12.53 1.86 13.73 2.18 ;
        RECT  11.13 4.22 13.53 4.54 ;
        POLYGON  12.15 2.18 5.52 2.18 5.52 2.34 5.20 2.34 5.20 1.86 12.15 1.86 ;
        POLYGON  12.15 3.90 10.77 3.90 10.77 4.54 10.45 4.54 10.45 3.58
                 12.15 3.58 ;
        RECT  2.96 1.22 10.77 1.54 ;
        POLYGON  8.61 3.90 5.68 3.90 5.68 3.58 8.12 3.58 8.12 2.50 8.44 2.50
                 8.44 3.58 8.61 3.58 ;
        POLYGON  7.76 3.26 6.02 3.26 6.02 2.94 7.44 2.94 7.44 2.50 7.76 2.50 ;
        POLYGON  4.72 4.36 4.40 4.36 4.40 3.90 2.96 3.90 2.96 3.58 4.72 3.58 ;
        POLYGON  4.06 2.18 0.18 2.18 0.18 1.76 0.50 1.76 0.50 1.86 4.06 1.86 ;
        RECT  1.58 4.22 3.98 4.54 ;
        RECT  1.58 1.22 2.58 1.54 ;
        POLYGON  2.58 3.90 0.50 3.90 0.50 4.54 0.18 4.54 0.18 3.58 2.58 3.58 ;
    END
END mux4_4

MACRO mux4_2
    CLASS CORE ;
    FOREIGN mux4_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 17.28 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  14.05 2.08 14.56 2.62 ;
        END
    END d0
    PIN d1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  14.88 1.98 15.20 2.62 ;
        END
    END d1
    PIN d2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.15 2.60 1.76 3.04 ;
        END
    END d2
    PIN d3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.60 0.83 3.04 ;
        END
    END d3
    PIN sl0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.80  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.26 2.50 3.68 3.04 ;
        END
    END sl0
    PIN sl1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.44 3.68 8.93 3.68 8.93 2.90 9.25 2.90 9.25 3.36 9.44 3.36 ;
        END
    END sl1
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  17.12 2.40 16.72 2.40 16.72 4.54 16.40 4.54 16.40 1.22
                 16.72 1.22 16.72 2.08 17.12 2.08 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 17.28 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  17.28 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 14.11 4.86 14.11 4.22 14.43 4.22 14.43 4.86
                 15.70 4.86 15.70 3.66 16.02 3.66 16.02 4.86 17.28 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  16.08 3.26 10.08 3.26 10.08 4.54 5.04 4.54 5.04 3.04 4.42 3.04
                 4.42 2.34 4.74 2.34 4.74 2.72 5.36 2.72 5.36 4.22 9.76 4.22
                 9.76 2.82 9.67 2.82 9.67 2.50 10.08 2.50 10.08 2.94 15.76 2.94
                 15.76 2.62 16.08 2.62 ;
        RECT  11.13 1.22 15.34 1.54 ;
        POLYGON  15.34 4.54 15.02 4.54 15.02 3.90 12.53 3.90 12.53 3.58
                 15.34 3.58 ;
        RECT  12.53 1.86 13.73 2.18 ;
        RECT  11.13 4.22 13.53 4.54 ;
        POLYGON  12.15 2.18 5.52 2.18 5.52 2.34 5.20 2.34 5.20 1.86 12.15 1.86 ;
        POLYGON  12.15 3.90 10.77 3.90 10.77 4.54 10.45 4.54 10.45 3.58
                 12.15 3.58 ;
        RECT  2.96 1.22 10.77 1.54 ;
        POLYGON  8.61 3.90 5.68 3.90 5.68 3.58 8.12 3.58 8.12 2.50 8.44 2.50
                 8.44 3.58 8.61 3.58 ;
        POLYGON  7.76 3.26 6.02 3.26 6.02 2.94 7.44 2.94 7.44 2.50 7.76 2.50 ;
        POLYGON  4.72 4.36 4.40 4.36 4.40 3.90 2.96 3.90 2.96 3.58 4.72 3.58 ;
        POLYGON  4.06 2.18 0.18 2.18 0.18 1.76 0.50 1.76 0.50 1.86 4.06 1.86 ;
        RECT  1.58 4.22 3.98 4.54 ;
        RECT  1.58 1.22 2.58 1.54 ;
        POLYGON  2.58 3.90 0.50 3.90 0.50 4.54 0.18 4.54 0.18 3.58 2.58 3.58 ;
    END
END mux4_2

MACRO mux4_1
    CLASS CORE ;
    FOREIGN mux4_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 17.28 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  14.05 2.08 14.56 2.62 ;
        END
    END d0
    PIN d1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  14.88 1.98 15.20 2.62 ;
        END
    END d1
    PIN d2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.15 2.60 1.76 3.04 ;
        END
    END d2
    PIN d3
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.60 0.83 3.04 ;
        END
    END d3
    PIN sl0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.80  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.26 2.50 3.68 3.04 ;
        END
    END sl0
    PIN sl1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.44 3.68 8.93 3.68 8.93 2.90 9.25 2.90 9.25 3.36 9.44 3.36 ;
        END
    END sl1
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  17.12 2.40 16.72 2.40 16.72 4.54 16.40 4.54 16.40 1.22
                 16.72 1.22 16.72 2.08 17.12 2.08 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 17.28 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  17.28 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 14.11 4.86 14.11 4.22 14.43 4.22 14.43 4.86
                 15.70 4.86 15.70 4.22 16.02 4.22 16.02 4.86 17.28 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  16.08 3.26 10.08 3.26 10.08 4.54 5.04 4.54 5.04 3.04 4.42 3.04
                 4.42 2.34 4.74 2.34 4.74 2.72 5.36 2.72 5.36 4.22 9.76 4.22
                 9.76 2.82 9.67 2.82 9.67 2.50 10.08 2.50 10.08 2.94 15.76 2.94
                 15.76 2.62 16.08 2.62 ;
        RECT  11.13 1.22 15.34 1.54 ;
        POLYGON  15.34 4.54 15.02 4.54 15.02 3.90 12.53 3.90 12.53 3.58
                 15.34 3.58 ;
        RECT  12.53 1.86 13.73 2.18 ;
        RECT  11.13 4.22 13.53 4.54 ;
        POLYGON  12.15 2.18 5.52 2.18 5.52 2.34 5.20 2.34 5.20 1.86 12.15 1.86 ;
        POLYGON  12.15 3.90 10.77 3.90 10.77 4.54 10.45 4.54 10.45 3.58
                 12.15 3.58 ;
        RECT  2.96 1.22 10.77 1.54 ;
        POLYGON  8.61 3.90 5.68 3.90 5.68 3.58 8.12 3.58 8.12 2.50 8.44 2.50
                 8.44 3.58 8.61 3.58 ;
        POLYGON  7.76 3.26 6.02 3.26 6.02 2.94 7.44 2.94 7.44 2.50 7.76 2.50 ;
        POLYGON  4.72 4.36 4.40 4.36 4.40 3.90 2.96 3.90 2.96 3.58 4.72 3.58 ;
        POLYGON  4.06 2.18 0.18 2.18 0.18 1.76 0.50 1.76 0.50 1.86 4.06 1.86 ;
        RECT  1.58 4.22 3.98 4.54 ;
        RECT  1.58 1.22 2.58 1.54 ;
        POLYGON  2.58 3.90 0.50 3.90 0.50 4.54 0.18 4.54 0.18 3.58 2.58 3.58 ;
    END
END mux4_1

MACRO mux2_4
    CLASS CORE ;
    FOREIGN mux2_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.96 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 1.98 5.60 2.62 ;
        END
    END d0
    PIN d1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.92 1.98 6.24 2.62 ;
        END
    END d1
    PIN sl0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.17  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.72 1.44 3.04 ;
        END
    END sl0
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.65 4.54 8.33 4.54 8.33 3.98 7.25 3.98 7.25 4.54 6.93 4.54
                 6.93 3.66 8.33 3.66 8.33 2.40 7.84 2.40 7.84 2.08 8.33 2.08
                 8.33 1.54 6.93 1.54 6.93 1.22 8.65 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.96 0.90 1.20 0.90 1.20 1.00 0.88 1.00 0.88 0.90 0.00 0.90
                 0.00 -0.90 8.96 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  8.96 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 5.34 4.86 5.34 4.22 5.66 4.22 5.66 4.86 7.63 4.86
                 7.63 4.30 7.95 4.30 7.95 4.86 8.96 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  7.31 3.26 3.38 3.26 3.38 3.42 3.06 3.42 3.06 2.18 2.39 2.18
                 2.39 1.86 3.38 1.86 3.38 2.94 6.99 2.94 6.99 2.62 7.31 2.62 ;
        RECT  1.56 1.22 6.57 1.54 ;
        POLYGON  6.57 4.54 6.25 4.54 6.25 3.90 3.76 3.90 3.76 3.58 6.57 3.58 ;
        RECT  3.76 1.86 4.96 2.18 ;
        RECT  1.56 4.22 4.76 4.54 ;
        POLYGON  2.74 3.90 0.50 3.90 0.50 4.06 0.16 4.06 0.16 1.44 0.50 1.44
                 0.50 1.76 0.48 1.76 0.48 3.58 2.42 3.58 2.42 2.62 2.74 2.62 ;
    END
END mux2_4

MACRO mux2_2
    CLASS CORE ;
    FOREIGN mux2_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.32 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 1.98 5.60 2.62 ;
        END
    END d0
    PIN d1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.92 1.98 6.24 2.62 ;
        END
    END d1
    PIN sl0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.17  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.72 1.44 3.04 ;
        END
    END sl0
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.16 2.40 7.95 2.40 7.95 4.54 7.63 4.54 7.63 1.22 7.95 1.22
                 7.95 2.08 8.16 2.08 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 0.90 7.25 0.90 7.25 1.54 6.93 1.54 6.93 0.90 1.20 0.90
                 1.20 1.00 0.88 1.00 0.88 0.90 0.00 0.90 0.00 -0.90 8.32 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 5.33 4.86 5.33 4.22 5.65 4.22 5.65 4.86 6.93 4.86
                 6.93 3.66 7.25 3.66 7.25 4.86 8.32 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  7.31 3.26 3.38 3.26 3.38 3.42 3.06 3.42 3.06 2.18 2.38 2.18
                 2.38 1.86 3.38 1.86 3.38 2.94 6.99 2.94 6.99 2.62 7.31 2.62 ;
        RECT  1.56 1.22 6.57 1.54 ;
        POLYGON  6.57 4.54 6.25 4.54 6.25 3.90 3.76 3.90 3.76 3.58 6.57 3.58 ;
        RECT  3.76 1.86 4.96 2.18 ;
        RECT  1.56 4.22 4.76 4.54 ;
        POLYGON  2.74 3.90 0.50 3.90 0.50 4.06 0.16 4.06 0.16 1.44 0.50 1.44
                 0.50 1.76 0.48 1.76 0.48 3.58 2.42 3.58 2.42 2.62 2.74 2.62 ;
    END
END mux2_2

MACRO mux2_1
    CLASS CORE ;
    FOREIGN mux2_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.32 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 1.98 5.60 2.62 ;
        END
    END d0
    PIN d1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.92 1.98 6.24 2.62 ;
        END
    END d1
    PIN sl0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.17  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.72 1.44 3.04 ;
        END
    END sl0
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.16 2.40 7.95 2.40 7.95 4.06 7.63 4.06 7.63 1.22 7.95 1.22
                 7.95 2.08 8.16 2.08 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 0.90 1.20 0.90 1.20 1.00 0.88 1.00 0.88 0.90 0.00 0.90
                 0.00 -0.90 8.32 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 5.34 4.86 5.34 4.22 5.66 4.22 5.66 4.86 6.93 4.86
                 6.93 4.14 7.25 4.14 7.25 4.86 8.32 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  7.31 3.26 3.38 3.26 3.38 3.42 3.06 3.42 3.06 2.18 2.39 2.18
                 2.39 1.86 3.38 1.86 3.38 2.94 7.31 2.94 ;
        RECT  1.56 1.22 6.57 1.54 ;
        POLYGON  6.57 4.46 6.25 4.46 6.25 3.90 3.76 3.90 3.76 3.58 6.57 3.58 ;
        RECT  3.76 1.86 4.96 2.18 ;
        RECT  1.56 4.22 4.76 4.54 ;
        POLYGON  2.74 3.90 0.50 3.90 0.50 4.06 0.16 4.06 0.16 1.44 0.50 1.44
                 0.50 1.76 0.48 1.76 0.48 3.58 2.42 3.58 2.42 2.62 2.74 2.62 ;
    END
END mux2_1

MACRO maj31_4
    CLASS CORE ;
    FOREIGN maj31_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 27.52 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        ANTENNAGATEAREA 1.14  LAYER metal2  ;
        ANTENNAMAXAREACAR 0.66  LAYER metal2  ;
        PORT
        LAYER metal2 ;
                POLYGON  22.66 2.40 2.96 2.40 2.96 3.04 2.64 3.04 2.64 2.08 22.66 2.08 ;
        LAYER v1 ;
        RECT  22.34 2.08 22.66 2.40 ;
        RECT  2.64 2.72 2.96 3.04 ;
        LAYER metal1 ;
        RECT  22.34 2.08 22.66 3.26 ;
        RECT  2.55 2.72 3.04 3.26 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.62 3.68 3.26 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        ANTENNAGATEAREA 1.14  LAYER metal2  ;
        ANTENNAMAXAREACAR 0.43  LAYER metal2  ;
        PORT
        LAYER metal2 ;
        RECT  4.64 2.72 22.02 3.04 ;
        LAYER v1 ;
        RECT  21.70 2.72 22.02 3.04 ;
        RECT  4.64 2.72 4.96 3.04 ;
        LAYER metal1 ;
        RECT  21.70 2.62 22.02 3.26 ;
        RECT  4.64 2.54 4.98 3.26 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.84  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  26.92 1.70 25.44 1.70 25.44 3.78 26.92 3.78 26.92 4.10
                 23.80 4.10 23.80 3.78 25.12 3.78 25.12 1.70 23.80 1.70
                 23.80 1.38 26.92 1.38 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 27.52 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 27.52 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  24.76 2.66 23.37 2.66 23.37 4.54 15.54 4.54 15.54 4.22
                 18.28 4.22 18.28 3.26 18.15 3.26 18.15 1.54 9.86 1.54
                 9.86 1.22 18.60 1.22 18.60 1.54 18.47 1.54 18.47 2.94
                 18.60 2.94 18.60 4.22 23.05 4.22 23.05 2.34 24.76 2.34 ;
        RECT  21.74 1.22 22.74 1.54 ;
        POLYGON  22.33 3.90 21.06 3.90 21.06 2.44 19.70 2.44 19.70 2.12
                 21.06 2.12 21.06 1.54 21.04 1.54 21.04 1.22 21.38 1.22
                 21.38 3.58 22.33 3.58 ;
        POLYGON  20.74 3.64 18.96 3.64 18.96 2.42 18.80 2.42 18.80 2.10
                 18.96 2.10 18.96 1.24 20.68 1.24 20.68 1.56 19.28 1.56
                 19.28 3.32 20.74 3.32 ;
        RECT  11.89 3.58 17.96 3.90 ;
        RECT  9.14 4.22 14.35 4.54 ;
        POLYGON  13.78 2.66 9.18 2.66 9.18 1.80 7.66 1.80 7.66 3.90 5.94 3.90
                 5.94 3.58 7.34 3.58 7.34 1.48 9.50 1.48 9.50 2.34 13.78 2.34 ;
        POLYGON  8.30 4.54 0.18 4.54 0.18 1.24 1.90 1.24 1.90 1.56 0.50 1.56
                 0.50 4.22 7.98 4.22 7.98 3.07 8.30 3.07 ;
        POLYGON  6.92 2.88 6.60 2.88 6.60 2.22 5.62 2.22 5.62 3.90 4.36 3.90
                 4.36 3.58 5.30 3.58 5.30 2.22 5.02 2.22 5.02 1.24 5.34 1.24
                 5.34 1.90 6.92 1.90 ;
        RECT  5.72 1.24 6.72 1.56 ;
        RECT  2.96 1.23 3.96 1.55 ;
        POLYGON  3.29 3.90 1.60 3.90 1.60 2.26 0.89 2.26 0.89 1.94 2.26 1.94
                 2.26 1.23 2.58 1.23 2.58 2.26 1.92 2.26 1.92 3.58 3.29 3.58 ;
    END
END maj31_4

MACRO maj31_2
    CLASS CORE ;
    FOREIGN maj31_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.84 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        ANTENNAGATEAREA 1.14  LAYER metal2  ;
        ANTENNAMAXAREACAR 0.66  LAYER metal2  ;
        PORT
        LAYER metal2 ;
                POLYGON  16.59 2.40 2.26 2.40 2.26 3.04 1.94 3.04 1.94 2.08 16.59 2.08 ;
        LAYER v1 ;
        RECT  16.27 2.08 16.59 2.40 ;
        RECT  1.94 2.72 2.26 3.04 ;
        LAYER metal1 ;
        RECT  16.27 2.08 16.59 3.26 ;
        RECT  1.85 2.72 2.40 3.26 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.62 3.04 3.26 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        ANTENNAGATEAREA 1.14  LAYER metal2  ;
        ANTENNAMAXAREACAR 0.40  LAYER metal2  ;
        PORT
        LAYER metal2 ;
        RECT  4.00 2.72 15.71 3.04 ;
        LAYER v1 ;
        RECT  15.39 2.72 15.71 3.04 ;
        RECT  4.00 2.72 4.32 3.04 ;
        LAYER metal1 ;
        RECT  15.39 2.62 15.71 3.26 ;
        RECT  4.00 2.54 4.32 3.26 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.04  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  19.68 4.54 17.49 4.54 17.49 4.22 19.36 4.22 19.36 1.70
                 17.49 1.70 17.49 1.38 19.68 1.38 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 19.84 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 19.84 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  18.45 2.66 17.23 2.66 17.23 3.90 17.17 3.90 17.17 4.54
                 11.80 4.54 11.80 4.22 13.14 4.22 13.14 3.26 12.55 3.26
                 12.55 1.54 9.16 1.54 9.16 1.22 12.87 1.22 12.87 2.94
                 13.46 2.94 13.46 4.22 16.85 4.22 16.85 3.58 16.91 3.58
                 16.91 2.34 18.45 2.34 ;
        POLYGON  16.46 3.90 14.75 3.90 14.75 2.44 14.52 2.44 14.52 2.12
                 14.75 2.12 14.75 1.54 14.73 1.54 14.73 1.22 15.07 1.22
                 15.07 3.58 16.46 3.58 ;
        RECT  15.43 1.22 16.43 1.54 ;
        POLYGON  14.20 3.64 13.88 3.64 13.88 2.42 13.19 2.42 13.19 2.10
                 13.35 2.10 13.35 1.24 13.67 1.24 13.67 2.10 14.20 2.10 ;
        RECT  9.71 3.58 12.82 3.90 ;
        POLYGON  10.87 2.66 8.48 2.66 8.48 1.82 6.66 1.82 6.66 3.90 5.94 3.90
                 5.94 3.58 6.34 3.58 6.34 1.50 8.80 1.50 8.80 2.34 10.87 2.34 ;
        RECT  8.31 4.22 10.75 4.54 ;
        POLYGON  7.50 4.54 0.18 4.54 0.18 1.24 0.50 1.24 0.50 4.22 7.18 4.22
                 7.18 3.07 7.50 3.07 ;
        RECT  5.02 1.24 6.02 1.56 ;
        POLYGON  5.96 2.86 4.96 2.86 4.96 3.90 3.66 3.90 3.66 3.58 4.64 3.58
                 4.64 2.22 4.32 2.22 4.32 1.24 4.64 1.24 4.64 1.90 4.96 1.90
                 4.96 2.54 5.96 2.54 ;
        RECT  2.26 1.23 3.26 1.55 ;
        POLYGON  2.59 3.90 0.90 3.90 0.90 2.26 0.89 2.26 0.89 1.94 1.56 1.94
                 1.56 1.23 1.88 1.23 1.88 2.26 1.22 2.26 1.22 3.58 2.59 3.58 ;
    END
END maj31_2

MACRO maj31_1
    CLASS CORE ;
    FOREIGN maj31_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.64 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        ANTENNAGATEAREA 1.14  LAYER metal2  ;
        ANTENNAMAXAREACAR 0.66  LAYER metal2  ;
        PORT
        LAYER metal2 ;
                POLYGON  14.63 2.40 2.26 2.40 2.26 3.04 1.94 3.04 1.94 2.08 14.63 2.08 ;
        LAYER v1 ;
        RECT  14.31 2.08 14.63 2.40 ;
        RECT  1.94 2.72 2.26 3.04 ;
        LAYER metal1 ;
        RECT  14.31 2.08 14.63 3.26 ;
        RECT  1.85 2.72 2.40 3.26 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.62 3.04 3.26 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        ANTENNAGATEAREA 1.14  LAYER metal2  ;
        ANTENNAMAXAREACAR 0.40  LAYER metal2  ;
        PORT
        LAYER metal2 ;
        RECT  4.00 2.72 13.75 3.04 ;
        LAYER v1 ;
        RECT  13.43 2.72 13.75 3.04 ;
        RECT  4.00 2.72 4.32 3.04 ;
        LAYER metal1 ;
        RECT  13.43 2.62 13.75 3.26 ;
        RECT  4.00 2.54 4.32 3.26 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.48 4.54 15.78 4.54 15.78 4.22 16.16 4.22 16.16 1.70
                 15.78 1.70 15.78 1.38 16.48 1.38 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 16.64 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 16.64 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  15.33 3.90 15.21 3.90 15.21 4.54 11.04 4.54 11.04 3.26
                 10.59 3.26 10.59 1.54 9.16 1.54 9.16 1.22 10.91 1.22
                 10.91 2.94 11.36 2.94 11.36 4.22 14.89 4.22 14.89 3.58
                 15.01 3.58 15.01 2.34 15.33 2.34 ;
        POLYGON  14.50 3.90 12.79 3.90 12.79 2.44 12.56 2.44 12.56 2.12
                 12.79 2.12 12.79 1.54 12.77 1.54 12.77 1.22 13.11 1.22
                 13.11 3.58 14.50 3.58 ;
        RECT  13.47 1.22 14.47 1.54 ;
        POLYGON  12.24 3.90 11.92 3.90 11.92 2.42 11.23 2.42 11.23 2.10
                 11.39 2.10 11.39 1.22 11.71 1.22 11.71 2.10 12.24 2.10 ;
        RECT  9.68 3.58 10.72 3.90 ;
        POLYGON  9.78 2.66 8.48 2.66 8.48 1.54 6.66 1.54 6.66 3.90 5.94 3.90
                 5.94 3.58 6.34 3.58 6.34 1.22 8.80 1.22 8.80 2.34 9.78 2.34 ;
        RECT  8.31 4.22 9.35 4.54 ;
        POLYGON  7.50 4.54 0.18 4.54 0.18 1.22 0.50 1.22 0.50 4.22 7.18 4.22
                 7.18 3.07 7.50 3.07 ;
        RECT  5.02 1.24 6.02 1.56 ;
        POLYGON  5.96 2.86 4.96 2.86 4.96 3.90 3.66 3.90 3.66 3.58 4.64 3.58
                 4.64 2.22 4.32 2.22 4.32 1.24 4.64 1.24 4.64 1.90 4.96 1.90
                 4.96 2.54 5.96 2.54 ;
        RECT  2.26 1.23 3.26 1.55 ;
        POLYGON  2.59 3.90 0.90 3.90 0.90 2.26 0.89 2.26 0.89 1.94 1.56 1.94
                 1.56 1.23 1.88 1.23 1.88 2.26 1.22 2.26 1.22 3.58 2.59 3.58 ;
    END
END maj31_1

MACRO latpsqb_4
    CLASS CORE ;
    FOREIGN latpsqb_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.64 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.00 2.02 11.32 2.02 11.32 1.70 11.68 1.70 11.68 1.44
                 12.00 1.44 ;
        END
    END gb
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.48 4.53 14.58 4.53 14.58 4.21 16.16 4.21 16.16 1.90
                 14.58 1.90 14.58 1.58 16.48 1.58 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.08 3.40 2.56 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 0.90 15.60 0.90 15.60 1.23 15.28 1.23 15.28 0.90
                 13.42 0.90 13.42 1.14 13.10 1.14 13.10 0.90 11.74 0.90
                 11.74 1.12 11.42 1.12 11.42 0.90 9.56 0.90 9.56 1.54 9.24 1.54
                 9.24 0.90 0.00 0.90 0.00 -0.90 16.64 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.82 2.58 4.82
                 2.58 4.86 2.94 4.86 2.94 4.62 3.26 4.62 3.26 4.86 9.34 4.86
                 9.34 4.16 9.66 4.16 9.66 4.86 11.42 4.86 11.42 4.16 11.74 4.16
                 11.74 4.86 16.64 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  15.60 3.89 13.08 3.89 13.08 4.54 12.76 4.54 12.76 3.89
                 12.32 3.89 12.32 1.22 12.64 1.22 12.64 3.57 15.28 3.57
                 15.28 2.34 15.60 2.34 ;
        POLYGON  14.12 1.90 14.10 1.90 14.10 3.08 13.78 3.08 13.78 1.58
                 14.12 1.58 ;
        POLYGON  11.90 2.68 11.68 2.68 11.68 3.84 8.79 3.84 8.79 3.90 6.77 3.90
                 6.77 3.84 5.42 3.84 5.42 4.30 5.10 4.30 5.10 1.22 5.42 1.22
                 5.42 3.52 7.09 3.52 7.09 3.58 8.47 3.58 8.47 3.52 11.36 3.52
                 11.36 2.36 11.90 2.36 ;
        POLYGON  11.04 1.54 11.00 1.54 11.00 2.88 11.04 2.88 11.04 3.20
                 10.68 3.20 10.68 2.48 10.56 2.48 10.56 2.16 10.68 2.16
                 10.68 1.22 11.04 1.22 ;
        POLYGON  10.36 3.20 9.92 3.20 9.92 2.44 6.47 2.44 6.47 2.12 9.92 2.12
                 9.92 1.22 10.26 1.22 10.26 1.54 10.24 1.54 10.24 2.88
                 10.36 2.88 ;
        POLYGON  8.98 4.54 5.80 4.54 5.80 4.16 6.12 4.16 6.12 4.22 8.98 4.22 ;
        RECT  5.80 1.22 8.86 1.54 ;
        RECT  7.28 2.94 8.28 3.26 ;
        RECT  0.18 1.22 4.72 1.54 ;
        POLYGON  4.72 4.30 2.50 4.30 2.50 4.50 0.50 4.50 0.50 4.54 0.18 4.54
                 0.18 4.18 2.18 4.18 2.18 3.98 4.72 3.98 ;
        POLYGON  4.04 3.66 3.72 3.66 3.72 3.20 1.96 3.20 1.96 2.88 3.72 2.88
                 3.72 1.86 4.04 1.86 ;
        RECT  0.88 3.54 1.88 3.86 ;
    END
END latpsqb_4

MACRO latpsqb_2
    CLASS CORE ;
    FOREIGN latpsqb_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.00 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.00 2.02 11.32 2.02 11.32 1.70 11.68 1.70 11.68 1.44
                 12.00 1.44 ;
        END
    END gb
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.12  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  15.84 2.40 15.72 2.40 15.72 4.54 15.40 4.54 15.40 1.22
                 15.72 1.22 15.72 2.08 15.84 2.08 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.08 3.40 2.56 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 0.90 13.42 0.90 13.42 1.14 13.10 1.14 13.10 0.90
                 11.74 0.90 11.74 1.12 11.42 1.12 11.42 0.90 9.56 0.90
                 9.56 1.54 9.24 1.54 9.24 0.90 0.00 0.90 0.00 -0.90 16.00 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.82 2.58 4.82
                 2.58 4.86 2.94 4.86 2.94 4.62 3.26 4.62 3.26 4.86 9.34 4.86
                 9.34 4.16 9.66 4.16 9.66 4.86 11.42 4.86 11.42 4.16 11.74 4.16
                 11.74 4.86 16.00 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  15.06 2.62 14.98 2.62 14.98 4.54 12.32 4.54 12.32 1.22
                 12.64 1.22 12.64 4.22 14.66 4.22 14.66 2.30 15.06 2.30 ;
        POLYGON  14.12 1.90 14.10 1.90 14.10 3.08 13.78 3.08 13.78 1.58
                 14.12 1.58 ;
        POLYGON  11.90 2.68 11.68 2.68 11.68 3.84 8.79 3.84 8.79 3.90 6.77 3.90
                 6.77 3.84 5.42 3.84 5.42 4.30 5.10 4.30 5.10 1.22 5.42 1.22
                 5.42 3.52 7.09 3.52 7.09 3.58 8.47 3.58 8.47 3.52 11.36 3.52
                 11.36 2.36 11.90 2.36 ;
        POLYGON  11.04 1.54 11.00 1.54 11.00 2.88 11.04 2.88 11.04 3.20
                 10.68 3.20 10.68 2.48 10.56 2.48 10.56 2.16 10.68 2.16
                 10.68 1.22 11.04 1.22 ;
        POLYGON  10.36 3.20 9.92 3.20 9.92 2.44 6.47 2.44 6.47 2.12 9.92 2.12
                 9.92 1.22 10.26 1.22 10.26 1.54 10.24 1.54 10.24 2.88
                 10.36 2.88 ;
        POLYGON  8.98 4.54 5.80 4.54 5.80 4.16 6.12 4.16 6.12 4.22 8.98 4.22 ;
        RECT  5.80 1.22 8.86 1.54 ;
        RECT  7.28 2.94 8.28 3.26 ;
        RECT  0.18 1.22 4.72 1.54 ;
        POLYGON  4.72 4.30 2.50 4.30 2.50 4.50 0.50 4.50 0.50 4.54 0.18 4.54
                 0.18 4.18 2.18 4.18 2.18 3.98 4.72 3.98 ;
        POLYGON  4.04 3.66 3.72 3.66 3.72 3.20 1.96 3.20 1.96 2.88 3.72 2.88
                 3.72 1.86 4.04 1.86 ;
        RECT  0.88 3.54 1.88 3.86 ;
    END
END latpsqb_2

MACRO latpsqb_1
    CLASS CORE ;
    FOREIGN latpsqb_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.00 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.00 2.02 11.32 2.02 11.32 1.70 11.68 1.70 11.68 1.44
                 12.00 1.44 ;
        END
    END gb
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  15.84 2.40 15.72 2.40 15.72 4.54 15.40 4.54 15.40 1.22
                 15.72 1.22 15.72 2.08 15.84 2.08 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.08 3.40 2.56 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 0.90 13.42 0.90 13.42 1.14 13.10 1.14 13.10 0.90
                 11.74 0.90 11.74 1.12 11.42 1.12 11.42 0.90 9.56 0.90
                 9.56 1.54 9.24 1.54 9.24 0.90 0.00 0.90 0.00 -0.90 16.00 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.82 2.58 4.82
                 2.58 4.86 2.94 4.86 2.94 4.62 3.26 4.62 3.26 4.86 9.34 4.86
                 9.34 4.16 9.66 4.16 9.66 4.86 11.42 4.86 11.42 4.16 11.74 4.16
                 11.74 4.86 16.00 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  15.06 2.62 14.98 2.62 14.98 4.54 12.32 4.54 12.32 1.22
                 12.64 1.22 12.64 4.22 14.66 4.22 14.66 2.30 15.06 2.30 ;
        POLYGON  14.12 1.90 14.10 1.90 14.10 3.08 13.78 3.08 13.78 1.58
                 14.12 1.58 ;
        POLYGON  11.90 2.68 11.68 2.68 11.68 3.84 8.79 3.84 8.79 3.90 6.77 3.90
                 6.77 3.84 5.42 3.84 5.42 4.30 5.10 4.30 5.10 1.22 5.42 1.22
                 5.42 3.52 7.09 3.52 7.09 3.58 8.47 3.58 8.47 3.52 11.36 3.52
                 11.36 2.36 11.90 2.36 ;
        POLYGON  11.04 1.54 11.00 1.54 11.00 2.88 11.04 2.88 11.04 3.20
                 10.68 3.20 10.68 2.48 10.56 2.48 10.56 2.16 10.68 2.16
                 10.68 1.22 11.04 1.22 ;
        POLYGON  10.36 3.20 9.92 3.20 9.92 2.44 6.47 2.44 6.47 2.12 9.92 2.12
                 9.92 1.22 10.26 1.22 10.26 1.54 10.24 1.54 10.24 2.88
                 10.36 2.88 ;
        POLYGON  8.98 4.54 5.80 4.54 5.80 4.16 6.12 4.16 6.12 4.22 8.98 4.22 ;
        RECT  5.80 1.22 8.86 1.54 ;
        RECT  7.28 2.94 8.28 3.26 ;
        RECT  0.18 1.22 4.72 1.54 ;
        POLYGON  4.72 4.30 2.50 4.30 2.50 4.50 0.50 4.50 0.50 4.54 0.18 4.54
                 0.18 4.18 2.18 4.18 2.18 3.98 4.72 3.98 ;
        POLYGON  4.04 3.66 3.72 3.66 3.72 3.20 1.96 3.20 1.96 2.88 3.72 2.88
                 3.72 1.86 4.04 1.86 ;
        RECT  0.88 3.54 1.88 3.86 ;
    END
END latpsqb_1

MACRO latpsq_4
    CLASS CORE ;
    FOREIGN latpsq_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.64 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.00 2.02 11.32 2.02 11.32 1.70 11.68 1.70 11.68 1.44
                 12.00 1.44 ;
        END
    END gb
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.48 3.25 13.99 3.25 13.99 2.93 16.16 2.93 16.16 1.62
                 14.48 1.62 14.48 1.30 16.48 1.30 ;
        END
    END q
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.08 3.40 2.56 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 0.90 13.42 0.90 13.42 1.14 13.10 1.14 13.10 0.90
                 11.74 0.90 11.74 1.12 11.42 1.12 11.42 0.90 9.56 0.90
                 9.56 1.54 9.24 1.54 9.24 0.90 0.00 0.90 0.00 -0.90 16.64 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.82 2.58 4.82
                 2.58 4.86 2.94 4.86 2.94 4.62 3.26 4.62 3.26 4.86 9.34 4.86
                 9.34 4.16 9.66 4.16 9.66 4.86 11.42 4.86 11.42 4.16 11.74 4.16
                 11.74 4.86 14.63 4.86 14.63 4.79 15.05 4.79 15.05 4.86
                 16.64 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  14.49 2.55 13.78 2.55 13.78 1.58 14.12 1.58 14.12 1.90
                 14.10 1.90 14.10 2.23 14.49 2.23 ;
        POLYGON  13.08 4.54 12.76 4.54 12.76 4.10 12.32 4.10 12.32 1.22
                 12.64 1.22 12.64 3.78 13.08 3.78 ;
        POLYGON  11.90 2.68 11.68 2.68 11.68 3.84 8.79 3.84 8.79 3.90 6.77 3.90
                 6.77 3.84 5.42 3.84 5.42 4.30 5.10 4.30 5.10 1.22 5.42 1.22
                 5.42 3.52 7.09 3.52 7.09 3.58 8.47 3.58 8.47 3.52 11.36 3.52
                 11.36 2.36 11.90 2.36 ;
        POLYGON  11.04 1.54 11.00 1.54 11.00 2.88 11.04 2.88 11.04 3.20
                 10.68 3.20 10.68 2.48 10.56 2.48 10.56 2.16 10.68 2.16
                 10.68 1.22 11.04 1.22 ;
        POLYGON  10.36 3.20 9.92 3.20 9.92 2.44 6.47 2.44 6.47 2.12 9.92 2.12
                 9.92 1.22 10.26 1.22 10.26 1.54 10.24 1.54 10.24 2.88
                 10.36 2.88 ;
        POLYGON  8.98 4.54 5.80 4.54 5.80 4.16 6.12 4.16 6.12 4.22 8.98 4.22 ;
        RECT  5.80 1.22 8.86 1.54 ;
        RECT  7.28 2.94 8.28 3.26 ;
        RECT  0.18 1.22 4.72 1.54 ;
        POLYGON  4.72 4.30 2.50 4.30 2.50 4.50 0.50 4.50 0.50 4.54 0.18 4.54
                 0.18 4.18 2.18 4.18 2.18 3.98 4.72 3.98 ;
        POLYGON  4.04 3.66 3.72 3.66 3.72 3.20 1.96 3.20 1.96 2.88 3.72 2.88
                 3.72 1.86 4.04 1.86 ;
        RECT  0.88 3.54 1.88 3.86 ;
    END
END latpsq_4

MACRO latpsq_2
    CLASS CORE ;
    FOREIGN latpsq_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.00 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.00 2.02 11.32 2.02 11.32 1.70 11.68 1.70 11.68 1.44
                 12.00 1.44 ;
        END
    END gb
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.80  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  15.20 1.76 14.76 1.76 14.76 4.54 14.42 4.54 14.42 3.14
                 14.44 3.14 14.44 1.22 14.80 1.22 14.80 1.44 15.20 1.44 ;
        END
    END q
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.08 3.40 2.56 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 0.90 13.42 0.90 13.42 1.14 13.10 1.14 13.10 0.90
                 11.74 0.90 11.74 1.12 11.42 1.12 11.42 0.90 9.56 0.90
                 9.56 1.54 9.24 1.54 9.24 0.90 0.00 0.90 0.00 -0.90 16.00 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.82 2.58 4.82
                 2.58 4.86 2.94 4.86 2.94 4.62 3.26 4.62 3.26 4.86 9.34 4.86
                 9.34 4.16 9.66 4.16 9.66 4.86 11.42 4.86 11.42 4.16 11.74 4.16
                 11.74 4.86 15.18 4.86 15.18 4.22 15.50 4.22 15.50 4.86
                 16.00 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  14.12 1.90 14.10 1.90 14.10 3.08 13.78 3.08 13.78 1.58
                 14.12 1.58 ;
        POLYGON  13.08 4.54 12.76 4.54 12.76 4.10 12.32 4.10 12.32 1.22
                 12.64 1.22 12.64 3.78 13.08 3.78 ;
        POLYGON  11.90 2.68 11.68 2.68 11.68 3.84 8.79 3.84 8.79 3.90 6.77 3.90
                 6.77 3.84 5.42 3.84 5.42 4.30 5.10 4.30 5.10 1.22 5.42 1.22
                 5.42 3.52 7.09 3.52 7.09 3.58 8.47 3.58 8.47 3.52 11.36 3.52
                 11.36 2.36 11.90 2.36 ;
        POLYGON  11.04 1.54 11.00 1.54 11.00 2.88 11.04 2.88 11.04 3.20
                 10.68 3.20 10.68 2.48 10.56 2.48 10.56 2.16 10.68 2.16
                 10.68 1.22 11.04 1.22 ;
        POLYGON  10.36 3.20 9.92 3.20 9.92 2.44 6.47 2.44 6.47 2.12 9.92 2.12
                 9.92 1.22 10.26 1.22 10.26 1.54 10.24 1.54 10.24 2.88
                 10.36 2.88 ;
        POLYGON  8.98 4.54 5.80 4.54 5.80 4.16 6.12 4.16 6.12 4.22 8.98 4.22 ;
        RECT  5.80 1.22 8.86 1.54 ;
        RECT  7.28 2.94 8.28 3.26 ;
        RECT  0.18 1.22 4.72 1.54 ;
        POLYGON  4.72 4.30 2.50 4.30 2.50 4.50 0.50 4.50 0.50 4.54 0.18 4.54
                 0.18 4.18 2.18 4.18 2.18 3.98 4.72 3.98 ;
        POLYGON  4.04 3.66 3.72 3.66 3.72 3.20 1.96 3.20 1.96 2.88 3.72 2.88
                 3.72 1.86 4.04 1.86 ;
        RECT  0.88 3.54 1.88 3.86 ;
    END
END latpsq_2

MACRO latpsq_1
    CLASS CORE ;
    FOREIGN latpsq_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.00 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.00 2.02 11.32 2.02 11.32 1.70 11.68 1.70 11.68 1.44
                 12.00 1.44 ;
        END
    END gb
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.29  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  15.20 1.76 14.76 1.76 14.76 4.54 14.44 4.54 14.44 1.22
                 14.80 1.22 14.80 1.44 15.20 1.44 ;
        END
    END q
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.08 3.40 2.56 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 0.90 13.42 0.90 13.42 1.14 13.10 1.14 13.10 0.90
                 11.74 0.90 11.74 1.12 11.42 1.12 11.42 0.90 9.56 0.90
                 9.56 1.54 9.24 1.54 9.24 0.90 0.00 0.90 0.00 -0.90 16.00 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.82 2.58 4.82
                 2.58 4.86 2.94 4.86 2.94 4.62 3.26 4.62 3.26 4.86 9.34 4.86
                 9.34 4.16 9.66 4.16 9.66 4.86 11.42 4.86 11.42 4.16 11.74 4.16
                 11.74 4.86 15.18 4.86 15.18 4.22 15.50 4.22 15.50 4.86
                 16.00 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  14.12 1.90 14.10 1.90 14.10 3.08 13.78 3.08 13.78 1.58
                 14.12 1.58 ;
        POLYGON  13.08 4.54 12.76 4.54 12.76 4.10 12.32 4.10 12.32 1.22
                 12.64 1.22 12.64 3.78 13.08 3.78 ;
        POLYGON  11.90 2.68 11.68 2.68 11.68 3.84 8.79 3.84 8.79 3.90 6.77 3.90
                 6.77 3.84 5.42 3.84 5.42 4.30 5.10 4.30 5.10 1.22 5.42 1.22
                 5.42 3.52 7.09 3.52 7.09 3.58 8.47 3.58 8.47 3.52 11.36 3.52
                 11.36 2.36 11.90 2.36 ;
        POLYGON  11.04 1.54 11.00 1.54 11.00 2.88 11.04 2.88 11.04 3.20
                 10.68 3.20 10.68 2.48 10.56 2.48 10.56 2.16 10.68 2.16
                 10.68 1.22 11.04 1.22 ;
        POLYGON  10.36 3.20 9.92 3.20 9.92 2.44 6.47 2.44 6.47 2.12 9.92 2.12
                 9.92 1.22 10.26 1.22 10.26 1.54 10.24 1.54 10.24 2.88
                 10.36 2.88 ;
        POLYGON  8.98 4.54 5.80 4.54 5.80 4.16 6.12 4.16 6.12 4.22 8.98 4.22 ;
        RECT  5.80 1.22 8.86 1.54 ;
        RECT  7.28 2.94 8.28 3.26 ;
        RECT  0.18 1.22 4.72 1.54 ;
        POLYGON  4.72 4.30 2.50 4.30 2.50 4.50 0.50 4.50 0.50 4.54 0.18 4.54
                 0.18 4.18 2.18 4.18 2.18 3.98 4.72 3.98 ;
        POLYGON  4.04 3.66 3.72 3.66 3.72 3.20 1.96 3.20 1.96 2.88 3.72 2.88
                 3.72 1.86 4.04 1.86 ;
        RECT  0.88 3.54 1.88 3.86 ;
    END
END latpsq_1

MACRO latps_4
    CLASS CORE ;
    FOREIGN latps_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.20 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.00 2.02 11.32 2.02 11.32 1.70 11.68 1.70 11.68 1.44
                 12.00 1.44 ;
        END
    END gb
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.73 3.25 14.96 3.25 14.96 2.93 16.16 2.93 16.16 2.72
                 16.41 2.72 16.41 1.62 14.48 1.62 14.48 1.30 16.73 1.30 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  19.04 4.53 17.05 4.53 17.05 4.21 18.72 4.21 18.72 1.90
                 17.05 1.90 17.05 1.58 19.04 1.58 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.08 3.40 2.56 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  19.20 0.90 18.07 0.90 18.07 1.23 17.75 1.23 17.75 0.90
                 13.42 0.90 13.42 1.14 13.10 1.14 13.10 0.90 11.74 0.90
                 11.74 1.12 11.42 1.12 11.42 0.90 9.56 0.90 9.56 1.54 9.24 1.54
                 9.24 0.90 0.00 0.90 0.00 -0.90 19.20 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  19.20 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.82 2.58 4.82
                 2.58 4.86 2.94 4.86 2.94 4.62 3.26 4.62 3.26 4.86 9.34 4.86
                 9.34 4.16 9.66 4.16 9.66 4.86 11.42 4.86 11.42 4.16 11.74 4.16
                 11.74 4.86 15.60 4.86 15.60 4.79 16.02 4.79 16.02 4.86
                 19.20 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  18.07 3.89 15.58 3.89 15.58 4.10 13.08 4.10 13.08 4.54
                 12.76 4.54 12.76 4.10 12.32 4.10 12.32 1.22 12.64 1.22
                 12.64 3.78 15.26 3.78 15.26 3.57 17.75 3.57 17.75 2.34
                 18.07 2.34 ;
        POLYGON  14.12 1.90 14.10 1.90 14.10 3.08 13.78 3.08 13.78 1.58
                 14.12 1.58 ;
        POLYGON  11.90 2.68 11.68 2.68 11.68 3.84 8.79 3.84 8.79 3.90 6.77 3.90
                 6.77 3.84 5.42 3.84 5.42 4.30 5.10 4.30 5.10 1.22 5.42 1.22
                 5.42 3.52 7.09 3.52 7.09 3.58 8.47 3.58 8.47 3.52 11.36 3.52
                 11.36 2.36 11.90 2.36 ;
        POLYGON  11.04 1.54 11.00 1.54 11.00 2.88 11.04 2.88 11.04 3.20
                 10.68 3.20 10.68 2.48 10.56 2.48 10.56 2.16 10.68 2.16
                 10.68 1.22 11.04 1.22 ;
        POLYGON  10.36 3.20 9.92 3.20 9.92 2.44 6.47 2.44 6.47 2.12 9.92 2.12
                 9.92 1.22 10.26 1.22 10.26 1.54 10.24 1.54 10.24 2.88
                 10.36 2.88 ;
        POLYGON  8.98 4.54 5.80 4.54 5.80 4.16 6.12 4.16 6.12 4.22 8.98 4.22 ;
        RECT  5.80 1.22 8.86 1.54 ;
        RECT  7.28 2.94 8.28 3.26 ;
        RECT  0.18 1.22 4.72 1.54 ;
        POLYGON  4.72 4.30 2.50 4.30 2.50 4.50 0.50 4.50 0.50 4.54 0.18 4.54
                 0.18 4.18 2.18 4.18 2.18 3.98 4.72 3.98 ;
        POLYGON  4.04 3.66 3.72 3.66 3.72 3.20 1.96 3.20 1.96 2.88 3.72 2.88
                 3.72 1.86 4.04 1.86 ;
        RECT  0.88 3.54 1.88 3.86 ;
    END
END latps_4

MACRO latps_2
    CLASS CORE ;
    FOREIGN latps_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.64 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.00 2.02 11.32 2.02 11.32 1.70 11.68 1.70 11.68 1.44
                 12.00 1.44 ;
        END
    END gb
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.84  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  15.20 1.76 14.76 1.76 14.76 3.80 14.40 3.80 14.40 3.48
                 14.44 3.48 14.44 1.22 14.80 1.22 14.80 1.44 15.20 1.44 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.12  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.48 2.40 16.32 2.40 16.32 4.54 16.00 4.54 16.00 1.22
                 16.32 1.22 16.32 2.08 16.48 2.08 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.08 3.40 2.56 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 0.90 13.42 0.90 13.42 1.14 13.10 1.14 13.10 0.90
                 11.74 0.90 11.74 1.12 11.42 1.12 11.42 0.90 9.56 0.90
                 9.56 1.54 9.24 1.54 9.24 0.90 0.00 0.90 0.00 -0.90 16.64 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.82 2.58 4.82
                 2.58 4.86 2.94 4.86 2.94 4.62 3.26 4.62 3.26 4.86 9.34 4.86
                 9.34 4.16 9.66 4.16 9.66 4.86 11.42 4.86 11.42 4.16 11.74 4.16
                 11.74 4.86 16.64 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  15.66 2.62 15.58 2.62 15.58 4.54 12.32 4.54 12.32 1.22
                 12.64 1.22 12.64 4.22 15.26 4.22 15.26 2.30 15.66 2.30 ;
        POLYGON  14.12 1.90 14.10 1.90 14.10 3.08 13.78 3.08 13.78 1.58
                 14.12 1.58 ;
        POLYGON  11.90 2.68 11.68 2.68 11.68 3.84 8.79 3.84 8.79 3.90 6.77 3.90
                 6.77 3.84 5.42 3.84 5.42 4.30 5.10 4.30 5.10 1.22 5.42 1.22
                 5.42 3.52 7.09 3.52 7.09 3.58 8.47 3.58 8.47 3.52 11.36 3.52
                 11.36 2.36 11.90 2.36 ;
        POLYGON  11.04 1.54 11.00 1.54 11.00 2.88 11.04 2.88 11.04 3.20
                 10.68 3.20 10.68 2.48 10.56 2.48 10.56 2.16 10.68 2.16
                 10.68 1.22 11.04 1.22 ;
        POLYGON  10.36 3.20 9.92 3.20 9.92 2.44 6.47 2.44 6.47 2.12 9.92 2.12
                 9.92 1.22 10.26 1.22 10.26 1.54 10.24 1.54 10.24 2.88
                 10.36 2.88 ;
        POLYGON  8.98 4.54 5.80 4.54 5.80 4.16 6.12 4.16 6.12 4.22 8.98 4.22 ;
        RECT  5.80 1.22 8.86 1.54 ;
        RECT  7.28 2.94 8.28 3.26 ;
        RECT  0.18 1.22 4.72 1.54 ;
        POLYGON  4.72 4.30 2.50 4.30 2.50 4.50 0.50 4.50 0.50 4.54 0.18 4.54
                 0.18 4.18 2.18 4.18 2.18 3.98 4.72 3.98 ;
        POLYGON  4.04 3.66 3.72 3.66 3.72 3.20 1.96 3.20 1.96 2.88 3.72 2.88
                 3.72 1.86 4.04 1.86 ;
        RECT  0.88 3.54 1.88 3.86 ;
    END
END latps_2

MACRO latps_1
    CLASS CORE ;
    FOREIGN latps_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.64 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.00 2.02 11.32 2.02 11.32 1.70 11.68 1.70 11.68 1.44
                 12.00 1.44 ;
        END
    END gb
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.43  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  15.20 1.76 14.76 1.76 14.76 3.65 14.40 3.65 14.40 3.33
                 14.44 3.33 14.44 1.22 14.80 1.22 14.80 1.44 15.20 1.44 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.48 2.40 16.32 2.40 16.32 4.54 16.00 4.54 16.00 1.22
                 16.32 1.22 16.32 2.08 16.48 2.08 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.08 3.40 2.56 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 0.90 13.42 0.90 13.42 1.14 13.10 1.14 13.10 0.90
                 11.74 0.90 11.74 1.12 11.42 1.12 11.42 0.90 9.56 0.90
                 9.56 1.54 9.24 1.54 9.24 0.90 0.00 0.90 0.00 -0.90 16.64 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.82 2.58 4.82
                 2.58 4.86 2.94 4.86 2.94 4.62 3.26 4.62 3.26 4.86 9.34 4.86
                 9.34 4.16 9.66 4.16 9.66 4.86 11.42 4.86 11.42 4.16 11.74 4.16
                 11.74 4.86 16.64 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  15.66 2.62 15.58 2.62 15.58 4.54 12.32 4.54 12.32 1.22
                 12.64 1.22 12.64 4.22 15.26 4.22 15.26 2.30 15.66 2.30 ;
        POLYGON  14.12 1.90 14.10 1.90 14.10 3.08 13.78 3.08 13.78 1.58
                 14.12 1.58 ;
        POLYGON  11.90 2.68 11.68 2.68 11.68 3.84 8.79 3.84 8.79 3.90 6.77 3.90
                 6.77 3.84 5.42 3.84 5.42 4.30 5.10 4.30 5.10 1.22 5.42 1.22
                 5.42 3.52 7.09 3.52 7.09 3.58 8.47 3.58 8.47 3.52 11.36 3.52
                 11.36 2.36 11.90 2.36 ;
        POLYGON  11.04 1.54 11.00 1.54 11.00 2.88 11.04 2.88 11.04 3.20
                 10.68 3.20 10.68 2.48 10.56 2.48 10.56 2.16 10.68 2.16
                 10.68 1.22 11.04 1.22 ;
        POLYGON  10.36 3.20 9.92 3.20 9.92 2.44 6.47 2.44 6.47 2.12 9.92 2.12
                 9.92 1.22 10.26 1.22 10.26 1.54 10.24 1.54 10.24 2.88
                 10.36 2.88 ;
        POLYGON  8.98 4.54 5.80 4.54 5.80 4.16 6.12 4.16 6.12 4.22 8.98 4.22 ;
        RECT  5.80 1.22 8.86 1.54 ;
        RECT  7.28 2.94 8.28 3.26 ;
        RECT  0.18 1.22 4.72 1.54 ;
        POLYGON  4.72 4.30 2.50 4.30 2.50 4.50 0.50 4.50 0.50 4.54 0.18 4.54
                 0.18 4.18 2.18 4.18 2.18 3.98 4.72 3.98 ;
        POLYGON  4.04 3.66 3.72 3.66 3.72 3.20 1.96 3.20 1.96 2.88 3.72 2.88
                 3.72 1.86 4.04 1.86 ;
        RECT  0.88 3.54 1.88 3.86 ;
    END
END latps_1

MACRO latprsqb_4
    CLASS CORE ;
    FOREIGN latprsqb_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.76 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.72 3.68 3.36 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.58 2.72 14.26 2.72 14.26 2.40 14.24 2.40 14.24 2.08
                 14.58 2.08 ;
        END
    END gb
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.37  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  21.60 2.40 21.23 2.40 21.23 4.54 19.38 4.54 19.38 4.22
                 20.91 4.22 20.91 1.54 19.39 1.54 19.39 1.22 21.23 1.22
                 21.23 2.08 21.60 2.08 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  18.08 1.22 18.59 1.86 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.90  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.71 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.76 0.90 17.69 0.90 17.69 1.28 17.37 1.28 17.37 0.90
                 14.78 0.90 14.78 1.14 14.46 1.14 14.46 0.90 12.60 0.90
                 12.60 1.28 12.28 1.28 12.28 0.90 8.24 0.90 8.24 1.24 7.92 1.24
                 7.92 0.90 1.20 0.90 1.20 1.28 0.88 1.28 0.88 0.90 0.00 0.90
                 0.00 -0.90 21.76 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.76 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.16 1.20 4.16
                 1.20 4.86 1.56 4.86 1.56 4.16 1.88 4.16 1.88 4.86 12.28 4.86
                 12.28 4.16 12.60 4.16 12.60 4.86 14.42 4.86 14.42 4.16
                 15.30 4.16 15.30 4.86 16.67 4.86 16.67 2.95 16.99 2.95
                 16.99 4.86 21.76 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.49 3.90 19.04 3.90 19.04 4.54 17.43 4.54 17.43 2.52
                 16.21 2.52 16.21 3.21 15.89 3.21 15.89 2.18 15.46 2.18
                 15.28 2.00 15.28 1.22 15.60 1.22 15.60 1.86 16.21 1.86
                 16.21 2.20 17.75 2.20 17.75 4.22 18.72 4.22 18.72 3.58
                 20.17 3.58 20.17 2.30 20.49 2.30 ;
        RECT  18.71 2.36 19.05 3.26 ;
        RECT  15.98 1.22 16.99 1.54 ;
        POLYGON  15.22 3.84 5.34 3.84 5.34 4.30 5.02 4.30 5.02 3.52 5.18 3.52
                 5.18 1.90 5.50 1.90 5.50 3.52 14.90 3.52 14.90 2.40 15.22 2.40 ;
        POLYGON  14.08 1.54 13.94 1.54 13.94 1.95 13.82 2.07 13.82 2.48
                 13.94 2.60 13.94 2.88 13.98 2.88 13.98 3.20 13.62 3.20
                 13.62 2.74 13.50 2.62 13.50 1.93 13.62 1.81 13.62 1.22
                 14.08 1.22 ;
        POLYGON  13.30 1.62 13.18 1.74 13.18 2.88 13.30 2.88 13.30 3.20
                 6.16 3.20 6.16 2.88 12.86 2.88 12.86 1.47 12.91 1.47
                 12.91 1.37 12.98 1.37 12.98 1.30 13.30 1.30 ;
        POLYGON  11.92 1.60 11.60 1.60 11.60 1.54 8.88 1.54 8.88 1.88 7.28 1.88
                 7.28 1.60 6.46 1.60 6.46 1.28 7.60 1.28 7.60 1.56 8.56 1.56
                 8.56 1.22 11.92 1.22 ;
        POLYGON  11.92 4.54 5.72 4.54 5.72 4.16 6.04 4.16 6.04 4.22 11.92 4.22 ;
        POLYGON  11.22 2.52 8.70 2.52 8.70 2.20 10.90 2.20 10.90 2.04
                 11.22 2.04 ;
        POLYGON  7.46 2.52 5.82 2.52 5.82 1.54 4.86 1.54 4.86 2.24 2.52 2.24
                 2.52 1.22 2.84 1.22 2.84 1.92 4.54 1.92 4.54 1.22 6.14 1.22
                 6.14 2.20 7.46 2.20 ;
        POLYGON  4.64 4.30 3.96 4.30 3.96 4.54 3.64 4.54 3.64 3.98 4.64 3.98 ;
        POLYGON  4.22 1.60 3.90 1.60 3.90 1.54 3.22 1.54 3.22 1.22 4.22 1.22 ;
        RECT  2.26 4.22 3.26 4.54 ;
        POLYGON  2.18 3.42 0.50 3.42 0.50 4.48 0.16 4.48 0.16 1.22 0.50 1.22
                 0.50 1.54 0.48 1.54 0.48 3.10 2.18 3.10 ;
    END
END latprsqb_4

MACRO latprsqb_2
    CLASS CORE ;
    FOREIGN latprsqb_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.72 3.68 3.36 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.58 2.72 14.26 2.72 14.26 2.40 14.24 2.40 14.24 2.08
                 14.58 2.08 ;
        END
    END gb
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.71  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.96 2.40 20.53 2.40 20.53 4.54 20.11 4.54 20.11 4.22
                 20.21 4.22 20.21 1.54 20.09 1.54 20.09 1.22 20.53 1.22
                 20.53 2.08 20.96 2.08 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  18.08 1.22 18.59 1.86 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.90  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.71 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 0.90 19.71 0.90 19.71 1.26 19.39 1.26 19.39 0.90
                 17.69 0.90 17.69 1.28 17.37 1.28 17.37 0.90 14.78 0.90
                 14.78 1.14 14.46 1.14 14.46 0.90 12.60 0.90 12.60 1.28
                 12.28 1.28 12.28 0.90 8.24 0.90 8.24 1.24 7.92 1.24 7.92 0.90
                 1.20 0.90 1.20 1.28 0.88 1.28 0.88 0.90 0.00 0.90 0.00 -0.90
                 21.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.16 1.20 4.16
                 1.20 4.86 1.56 4.86 1.56 4.16 1.88 4.16 1.88 4.86 12.28 4.86
                 12.28 4.16 12.60 4.16 12.60 4.86 14.42 4.86 14.42 4.16
                 15.30 4.16 15.30 4.86 16.67 4.86 16.67 2.95 16.99 2.95
                 16.99 4.86 21.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  19.87 2.62 19.79 2.62 19.79 4.54 17.43 4.54 17.43 2.52
                 16.21 2.52 16.21 3.21 15.89 3.21 15.89 2.18 15.46 2.18
                 15.28 2.00 15.28 1.22 15.60 1.22 15.60 1.86 16.21 1.86
                 16.21 2.20 17.75 2.20 17.75 4.22 19.47 4.22 19.47 2.30
                 19.87 2.30 ;
        RECT  18.71 2.76 19.05 3.90 ;
        RECT  15.98 1.22 16.99 1.54 ;
        POLYGON  15.22 3.84 5.34 3.84 5.34 4.30 5.02 4.30 5.02 3.52 5.18 3.52
                 5.18 1.90 5.50 1.90 5.50 3.52 14.90 3.52 14.90 2.40 15.22 2.40 ;
        POLYGON  14.08 1.54 13.94 1.54 13.94 1.95 13.82 2.07 13.82 2.48
                 13.94 2.60 13.94 2.88 13.98 2.88 13.98 3.20 13.62 3.20
                 13.62 2.74 13.50 2.62 13.50 1.93 13.62 1.81 13.62 1.22
                 14.08 1.22 ;
        POLYGON  13.30 1.62 13.18 1.74 13.18 2.88 13.30 2.88 13.30 3.20
                 6.16 3.20 6.16 2.88 12.86 2.88 12.86 1.47 12.91 1.47
                 12.91 1.37 12.98 1.37 12.98 1.30 13.30 1.30 ;
        POLYGON  11.92 1.60 11.60 1.60 11.60 1.54 8.88 1.54 8.88 1.88 7.28 1.88
                 7.28 1.60 6.46 1.60 6.46 1.28 7.60 1.28 7.60 1.56 8.56 1.56
                 8.56 1.22 11.92 1.22 ;
        POLYGON  11.92 4.54 5.72 4.54 5.72 4.16 6.04 4.16 6.04 4.22 11.92 4.22 ;
        POLYGON  11.22 2.52 8.70 2.52 8.70 2.20 10.90 2.20 10.90 2.04
                 11.22 2.04 ;
        POLYGON  7.46 2.52 5.82 2.52 5.82 1.54 4.86 1.54 4.86 2.24 2.52 2.24
                 2.52 1.22 2.84 1.22 2.84 1.92 4.54 1.92 4.54 1.22 6.14 1.22
                 6.14 2.20 7.46 2.20 ;
        POLYGON  4.64 4.30 3.96 4.30 3.96 4.54 3.64 4.54 3.64 3.98 4.64 3.98 ;
        POLYGON  4.22 1.60 3.90 1.60 3.90 1.54 3.22 1.54 3.22 1.22 4.22 1.22 ;
        RECT  2.26 4.22 3.26 4.54 ;
        POLYGON  2.18 3.42 0.50 3.42 0.50 4.48 0.16 4.48 0.16 1.22 0.50 1.22
                 0.50 1.54 0.48 1.54 0.48 3.10 2.18 3.10 ;
    END
END latprsqb_2

MACRO latprsqb_1
    CLASS CORE ;
    FOREIGN latprsqb_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.72 3.68 3.36 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.58 2.72 14.26 2.72 14.26 2.40 14.24 2.40 14.24 2.08
                 14.58 2.08 ;
        END
    END gb
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.23  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.96 2.40 20.53 2.40 20.53 4.54 20.11 4.54 20.11 4.22
                 20.21 4.22 20.21 1.54 20.09 1.54 20.09 1.22 20.53 1.22
                 20.53 2.08 20.96 2.08 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  18.08 1.22 18.59 1.86 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.90  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.71 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 0.90 19.71 0.90 19.71 1.26 19.39 1.26 19.39 0.90
                 17.69 0.90 17.69 1.28 17.37 1.28 17.37 0.90 14.78 0.90
                 14.78 1.14 14.46 1.14 14.46 0.90 12.60 0.90 12.60 1.28
                 12.28 1.28 12.28 0.90 8.24 0.90 8.24 1.24 7.92 1.24 7.92 0.90
                 1.20 0.90 1.20 1.28 0.88 1.28 0.88 0.90 0.00 0.90 0.00 -0.90
                 21.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.16 1.20 4.16
                 1.20 4.86 1.56 4.86 1.56 4.16 1.88 4.16 1.88 4.86 12.28 4.86
                 12.28 4.16 12.60 4.16 12.60 4.86 14.42 4.86 14.42 4.16
                 15.30 4.16 15.30 4.86 16.67 4.86 16.67 2.95 16.99 2.95
                 16.99 4.86 21.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  19.87 2.62 19.79 2.62 19.79 4.54 17.43 4.54 17.43 2.52
                 16.21 2.52 16.21 3.21 15.89 3.21 15.89 2.18 15.46 2.18
                 15.28 2.00 15.28 1.22 15.60 1.22 15.60 1.86 16.21 1.86
                 16.21 2.20 17.75 2.20 17.75 4.22 19.47 4.22 19.47 2.30
                 19.87 2.30 ;
        RECT  18.71 2.76 19.05 3.90 ;
        RECT  15.98 1.22 16.99 1.54 ;
        POLYGON  15.22 3.84 5.34 3.84 5.34 4.30 5.02 4.30 5.02 3.52 5.18 3.52
                 5.18 1.90 5.50 1.90 5.50 3.52 14.90 3.52 14.90 2.40 15.22 2.40 ;
        POLYGON  14.08 1.54 13.94 1.54 13.94 1.95 13.82 2.07 13.82 2.48
                 13.94 2.60 13.94 2.88 13.98 2.88 13.98 3.20 13.62 3.20
                 13.62 2.74 13.50 2.62 13.50 1.93 13.62 1.81 13.62 1.22
                 14.08 1.22 ;
        POLYGON  13.30 1.62 13.18 1.74 13.18 2.88 13.30 2.88 13.30 3.20
                 6.16 3.20 6.16 2.88 12.86 2.88 12.86 1.47 12.91 1.47
                 12.91 1.37 12.98 1.37 12.98 1.30 13.30 1.30 ;
        POLYGON  11.92 1.60 11.60 1.60 11.60 1.54 8.88 1.54 8.88 1.88 7.28 1.88
                 7.28 1.60 6.46 1.60 6.46 1.28 7.60 1.28 7.60 1.56 8.56 1.56
                 8.56 1.22 11.92 1.22 ;
        POLYGON  11.92 4.54 5.72 4.54 5.72 4.16 6.04 4.16 6.04 4.22 11.92 4.22 ;
        POLYGON  11.22 2.52 8.70 2.52 8.70 2.20 10.90 2.20 10.90 2.04
                 11.22 2.04 ;
        POLYGON  7.46 2.52 5.82 2.52 5.82 1.54 4.86 1.54 4.86 2.24 2.52 2.24
                 2.52 1.22 2.84 1.22 2.84 1.92 4.54 1.92 4.54 1.22 6.14 1.22
                 6.14 2.20 7.46 2.20 ;
        POLYGON  4.64 4.30 3.96 4.30 3.96 4.54 3.64 4.54 3.64 3.98 4.64 3.98 ;
        POLYGON  4.22 1.60 3.90 1.60 3.90 1.54 3.22 1.54 3.22 1.22 4.22 1.22 ;
        RECT  2.26 4.22 3.26 4.54 ;
        POLYGON  2.18 3.42 0.50 3.42 0.50 4.48 0.16 4.48 0.16 1.22 0.50 1.22
                 0.50 1.54 0.48 1.54 0.48 3.10 2.18 3.10 ;
    END
END latprsqb_1

MACRO latprsq_4
    CLASS CORE ;
    FOREIGN latprsq_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.76 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.72 3.68 3.36 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.58 2.72 14.26 2.72 14.26 2.40 14.24 2.40 14.24 2.08
                 14.58 2.08 ;
        END
    END gb
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  21.42 3.25 19.65 3.25 19.65 2.93 20.64 2.93 20.64 2.72
                 21.10 2.72 21.10 1.62 19.17 1.62 19.17 1.30 21.42 1.30 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  18.08 1.22 18.59 1.86 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.90  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.71 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.76 0.90 17.69 0.90 17.69 1.28 17.37 1.28 17.37 0.90
                 14.78 0.90 14.78 1.14 14.46 1.14 14.46 0.90 12.60 0.90
                 12.60 1.28 12.28 1.28 12.28 0.90 8.24 0.90 8.24 1.24 7.92 1.24
                 7.92 0.90 1.20 0.90 1.20 1.28 0.88 1.28 0.88 0.90 0.00 0.90
                 0.00 -0.90 21.76 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.76 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.16 1.20 4.16
                 1.20 4.86 1.56 4.86 1.56 4.16 1.88 4.16 1.88 4.86 12.28 4.86
                 12.28 4.16 12.60 4.16 12.60 4.86 14.42 4.86 14.42 4.16
                 15.30 4.16 15.30 4.86 16.67 4.86 16.67 2.95 16.99 2.95
                 16.99 4.86 20.29 4.86 20.29 4.79 20.71 4.79 20.71 4.86
                 21.76 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  18.73 2.23 19.05 3.90 ;
        POLYGON  17.75 4.54 17.43 4.54 17.43 2.52 16.21 2.52 16.21 3.21
                 15.89 3.21 15.89 2.18 15.46 2.18 15.28 2.00 15.28 1.22
                 15.60 1.22 15.60 1.86 16.21 1.86 16.21 2.20 17.75 2.20 ;
        RECT  15.98 1.22 16.99 1.54 ;
        POLYGON  15.22 3.84 5.34 3.84 5.34 4.30 5.02 4.30 5.02 3.52 5.18 3.52
                 5.18 1.90 5.50 1.90 5.50 3.52 14.90 3.52 14.90 2.40 15.22 2.40 ;
        POLYGON  14.08 1.54 13.94 1.54 13.94 1.95 13.82 2.07 13.82 2.48
                 13.94 2.60 13.94 2.88 13.98 2.88 13.98 3.20 13.62 3.20
                 13.62 2.74 13.50 2.62 13.50 1.93 13.62 1.81 13.62 1.22
                 14.08 1.22 ;
        POLYGON  13.30 1.62 13.18 1.74 13.18 2.88 13.30 2.88 13.30 3.20
                 6.16 3.20 6.16 2.88 12.86 2.88 12.86 1.47 12.91 1.47
                 12.91 1.37 12.98 1.37 12.98 1.30 13.30 1.30 ;
        POLYGON  11.92 1.60 11.60 1.60 11.60 1.54 8.88 1.54 8.88 1.88 7.28 1.88
                 7.28 1.60 6.46 1.60 6.46 1.28 7.60 1.28 7.60 1.56 8.56 1.56
                 8.56 1.22 11.92 1.22 ;
        POLYGON  11.92 4.54 5.72 4.54 5.72 4.16 6.04 4.16 6.04 4.22 11.92 4.22 ;
        POLYGON  11.22 2.52 8.70 2.52 8.70 2.20 10.90 2.20 10.90 2.04
                 11.22 2.04 ;
        POLYGON  7.46 2.52 5.82 2.52 5.82 1.54 4.86 1.54 4.86 2.24 2.52 2.24
                 2.52 1.22 2.84 1.22 2.84 1.92 4.54 1.92 4.54 1.22 6.14 1.22
                 6.14 2.20 7.46 2.20 ;
        POLYGON  4.64 4.30 3.96 4.30 3.96 4.54 3.64 4.54 3.64 3.98 4.64 3.98 ;
        POLYGON  4.22 1.60 3.90 1.60 3.90 1.54 3.22 1.54 3.22 1.22 4.22 1.22 ;
        RECT  2.26 4.22 3.26 4.54 ;
        POLYGON  2.18 3.42 0.50 3.42 0.50 4.48 0.16 4.48 0.16 1.22 0.50 1.22
                 0.50 1.54 0.48 1.54 0.48 3.10 2.18 3.10 ;
    END
END latprsq_4

MACRO latprsq_2
    CLASS CORE ;
    FOREIGN latprsq_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 20.48 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.72 3.68 3.36 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.58 2.72 14.26 2.72 14.26 2.40 14.24 2.40 14.24 2.08
                 14.58 2.08 ;
        END
    END gb
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.32 1.76 20.27 1.76 20.27 4.54 19.95 4.54 19.95 1.22
                 20.27 1.22 20.27 1.44 20.32 1.44 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  18.08 1.22 18.59 1.86 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.90  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.71 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 0.90 19.57 0.90 19.57 1.26 19.25 1.26 19.25 0.90
                 17.69 0.90 17.69 1.28 17.37 1.28 17.37 0.90 14.78 0.90
                 14.78 1.14 14.46 1.14 14.46 0.90 12.60 0.90 12.60 1.28
                 12.28 1.28 12.28 0.90 8.24 0.90 8.24 1.24 7.92 1.24 7.92 0.90
                 1.20 0.90 1.20 1.28 0.88 1.28 0.88 0.90 0.00 0.90 0.00 -0.90
                 20.48 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.16 1.20 4.16
                 1.20 4.86 1.56 4.86 1.56 4.16 1.88 4.16 1.88 4.86 12.28 4.86
                 12.28 4.16 12.60 4.16 12.60 4.86 14.42 4.86 14.42 4.16
                 15.30 4.16 15.30 4.86 16.67 4.86 16.67 2.95 16.99 2.95
                 16.99 4.86 19.25 4.86 19.25 4.22 19.57 4.22 19.57 4.86
                 20.48 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  19.05 3.08 18.89 3.08 18.89 4.54 18.57 4.54 18.57 2.76
                 19.05 2.76 ;
        POLYGON  17.75 4.54 17.43 4.54 17.43 2.52 16.21 2.52 16.21 3.21
                 15.89 3.21 15.89 2.18 15.46 2.18 15.28 2.00 15.28 1.22
                 15.60 1.22 15.60 1.86 16.21 1.86 16.21 2.20 17.75 2.20 ;
        RECT  15.98 1.22 16.99 1.54 ;
        POLYGON  15.22 3.84 5.34 3.84 5.34 4.30 5.02 4.30 5.02 3.52 5.18 3.52
                 5.18 1.90 5.50 1.90 5.50 3.52 14.90 3.52 14.90 2.40 15.22 2.40 ;
        POLYGON  14.08 1.54 13.94 1.54 13.94 1.95 13.82 2.07 13.82 2.48
                 13.94 2.60 13.94 2.88 13.98 2.88 13.98 3.20 13.62 3.20
                 13.62 2.74 13.50 2.62 13.50 1.93 13.62 1.81 13.62 1.22
                 14.08 1.22 ;
        POLYGON  13.30 1.62 13.18 1.74 13.18 2.88 13.30 2.88 13.30 3.20
                 6.16 3.20 6.16 2.88 12.86 2.88 12.86 1.47 12.91 1.47
                 12.91 1.37 12.98 1.37 12.98 1.30 13.30 1.30 ;
        POLYGON  11.92 1.60 11.60 1.60 11.60 1.54 8.88 1.54 8.88 1.88 7.28 1.88
                 7.28 1.60 6.46 1.60 6.46 1.28 7.60 1.28 7.60 1.56 8.56 1.56
                 8.56 1.22 11.92 1.22 ;
        POLYGON  11.92 4.54 5.72 4.54 5.72 4.16 6.04 4.16 6.04 4.22 11.92 4.22 ;
        POLYGON  11.22 2.52 8.70 2.52 8.70 2.20 10.90 2.20 10.90 2.04
                 11.22 2.04 ;
        POLYGON  7.46 2.52 5.82 2.52 5.82 1.54 4.86 1.54 4.86 2.24 2.52 2.24
                 2.52 1.22 2.84 1.22 2.84 1.92 4.54 1.92 4.54 1.22 6.14 1.22
                 6.14 2.20 7.46 2.20 ;
        POLYGON  4.64 4.30 3.96 4.30 3.96 4.54 3.64 4.54 3.64 3.98 4.64 3.98 ;
        POLYGON  4.22 1.60 3.90 1.60 3.90 1.54 3.22 1.54 3.22 1.22 4.22 1.22 ;
        RECT  2.26 4.22 3.26 4.54 ;
        POLYGON  2.18 3.42 0.50 3.42 0.50 4.48 0.16 4.48 0.16 1.22 0.50 1.22
                 0.50 1.54 0.48 1.54 0.48 3.10 2.18 3.10 ;
    END
END latprsq_2

MACRO latprsq_1
    CLASS CORE ;
    FOREIGN latprsq_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 20.48 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.72 3.68 3.36 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.58 2.72 14.26 2.72 14.26 2.40 14.24 2.40 14.24 2.08
                 14.58 2.08 ;
        END
    END gb
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.32 1.76 20.27 1.76 20.27 4.54 19.95 4.54 19.95 1.22
                 20.27 1.22 20.27 1.44 20.32 1.44 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  18.08 1.22 18.59 1.86 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.90  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.71 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 0.90 19.57 0.90 19.57 1.26 19.25 1.26 19.25 0.90
                 17.69 0.90 17.69 1.28 17.37 1.28 17.37 0.90 14.78 0.90
                 14.78 1.14 14.46 1.14 14.46 0.90 12.60 0.90 12.60 1.28
                 12.28 1.28 12.28 0.90 8.24 0.90 8.24 1.24 7.92 1.24 7.92 0.90
                 1.20 0.90 1.20 1.28 0.88 1.28 0.88 0.90 0.00 0.90 0.00 -0.90
                 20.48 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.16 1.20 4.16
                 1.20 4.86 1.56 4.86 1.56 4.16 1.88 4.16 1.88 4.86 12.28 4.86
                 12.28 4.16 12.60 4.16 12.60 4.86 14.42 4.86 14.42 4.16
                 15.30 4.16 15.30 4.86 16.67 4.86 16.67 2.95 16.99 2.95
                 16.99 4.86 19.25 4.86 19.25 4.22 19.57 4.22 19.57 4.86
                 20.48 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  19.05 3.08 18.89 3.08 18.89 4.54 18.57 4.54 18.57 2.76
                 19.05 2.76 ;
        POLYGON  17.75 4.54 17.43 4.54 17.43 2.52 16.21 2.52 16.21 3.21
                 15.89 3.21 15.89 2.18 15.46 2.18 15.28 2.00 15.28 1.22
                 15.60 1.22 15.60 1.86 16.21 1.86 16.21 2.20 17.75 2.20 ;
        RECT  15.98 1.22 16.99 1.54 ;
        POLYGON  15.22 3.84 5.34 3.84 5.34 4.30 5.02 4.30 5.02 3.52 5.18 3.52
                 5.18 1.90 5.50 1.90 5.50 3.52 14.90 3.52 14.90 2.40 15.22 2.40 ;
        POLYGON  14.08 1.54 13.94 1.54 13.94 1.95 13.82 2.07 13.82 2.48
                 13.94 2.60 13.94 2.88 13.98 2.88 13.98 3.20 13.62 3.20
                 13.62 2.74 13.50 2.62 13.50 1.93 13.62 1.81 13.62 1.22
                 14.08 1.22 ;
        POLYGON  13.30 1.62 13.18 1.74 13.18 2.88 13.30 2.88 13.30 3.20
                 6.16 3.20 6.16 2.88 12.86 2.88 12.86 1.47 12.91 1.47
                 12.91 1.37 12.98 1.37 12.98 1.30 13.30 1.30 ;
        POLYGON  11.92 1.60 11.60 1.60 11.60 1.54 8.88 1.54 8.88 1.88 7.28 1.88
                 7.28 1.60 6.46 1.60 6.46 1.28 7.60 1.28 7.60 1.56 8.56 1.56
                 8.56 1.22 11.92 1.22 ;
        POLYGON  11.92 4.54 5.72 4.54 5.72 4.16 6.04 4.16 6.04 4.22 11.92 4.22 ;
        POLYGON  11.22 2.52 8.70 2.52 8.70 2.20 10.90 2.20 10.90 2.04
                 11.22 2.04 ;
        POLYGON  7.46 2.52 5.82 2.52 5.82 1.54 4.86 1.54 4.86 2.24 2.52 2.24
                 2.52 1.22 2.84 1.22 2.84 1.92 4.54 1.92 4.54 1.22 6.14 1.22
                 6.14 2.20 7.46 2.20 ;
        POLYGON  4.64 4.30 3.96 4.30 3.96 4.54 3.64 4.54 3.64 3.98 4.64 3.98 ;
        POLYGON  4.22 1.60 3.90 1.60 3.90 1.54 3.22 1.54 3.22 1.22 4.22 1.22 ;
        RECT  2.26 4.22 3.26 4.54 ;
        POLYGON  2.18 3.42 0.50 3.42 0.50 4.48 0.16 4.48 0.16 1.22 0.50 1.22
                 0.50 1.54 0.48 1.54 0.48 3.10 2.18 3.10 ;
    END
END latprsq_1

MACRO latprs_4
    CLASS CORE ;
    FOREIGN latprs_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.72 3.68 3.36 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.58 2.72 14.26 2.72 14.26 2.40 14.24 2.40 14.24 2.08
                 14.58 2.08 ;
        END
    END gb
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  21.42 3.25 19.65 3.25 19.65 2.93 20.64 2.93 20.64 2.72
                 21.10 2.72 21.10 1.62 19.17 1.62 19.17 1.30 21.42 1.30 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  23.52 4.53 21.74 4.53 21.74 4.21 23.20 4.21 23.20 1.90
                 21.74 1.90 21.74 1.58 23.52 1.58 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  18.08 1.22 18.59 1.86 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.90  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.71 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  23.68 0.90 22.76 0.90 22.76 1.23 22.44 1.23 22.44 0.90
                 17.69 0.90 17.69 1.28 17.37 1.28 17.37 0.90 14.78 0.90
                 14.78 1.14 14.46 1.14 14.46 0.90 12.60 0.90 12.60 1.28
                 12.28 1.28 12.28 0.90 8.24 0.90 8.24 1.24 7.92 1.24 7.92 0.90
                 1.20 0.90 1.20 1.28 0.88 1.28 0.88 0.90 0.00 0.90 0.00 -0.90
                 23.68 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  23.68 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.16 1.20 4.16
                 1.20 4.86 1.56 4.86 1.56 4.16 1.88 4.16 1.88 4.86 12.28 4.86
                 12.28 4.16 12.60 4.16 12.60 4.86 14.42 4.86 14.42 4.16
                 15.30 4.16 15.30 4.86 16.67 4.86 16.67 2.95 16.99 2.95
                 16.99 4.86 20.29 4.86 20.29 4.79 20.71 4.79 20.71 4.86
                 23.68 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  22.76 3.89 19.85 3.89 19.85 4.54 17.43 4.54 17.43 2.52
                 16.21 2.52 16.21 3.21 15.89 3.21 15.89 2.18 15.46 2.18
                 15.28 2.00 15.28 1.22 15.60 1.22 15.60 1.86 16.21 1.86
                 16.21 2.20 17.75 2.20 17.75 4.22 19.53 4.22 19.53 3.57
                 22.44 3.57 22.44 2.34 22.76 2.34 ;
        RECT  18.73 2.23 19.05 3.90 ;
        RECT  15.98 1.22 16.99 1.54 ;
        POLYGON  15.22 3.84 5.34 3.84 5.34 4.30 5.02 4.30 5.02 3.52 5.18 3.52
                 5.18 1.90 5.50 1.90 5.50 3.52 14.90 3.52 14.90 2.40 15.22 2.40 ;
        POLYGON  14.08 1.54 13.94 1.54 13.94 1.95 13.82 2.07 13.82 2.48
                 13.94 2.60 13.94 2.88 13.98 2.88 13.98 3.20 13.62 3.20
                 13.62 2.74 13.50 2.62 13.50 1.93 13.62 1.81 13.62 1.22
                 14.08 1.22 ;
        POLYGON  13.30 1.62 13.18 1.74 13.18 2.88 13.30 2.88 13.30 3.20
                 6.16 3.20 6.16 2.88 12.86 2.88 12.86 1.47 12.91 1.47
                 12.91 1.37 12.98 1.37 12.98 1.30 13.30 1.30 ;
        POLYGON  11.92 1.60 11.60 1.60 11.60 1.54 8.88 1.54 8.88 1.88 7.28 1.88
                 7.28 1.60 6.46 1.60 6.46 1.28 7.60 1.28 7.60 1.56 8.56 1.56
                 8.56 1.22 11.92 1.22 ;
        POLYGON  11.92 4.54 5.72 4.54 5.72 4.16 6.04 4.16 6.04 4.22 11.92 4.22 ;
        POLYGON  11.22 2.52 8.70 2.52 8.70 2.20 10.90 2.20 10.90 2.04
                 11.22 2.04 ;
        POLYGON  7.46 2.52 5.82 2.52 5.82 1.54 4.86 1.54 4.86 2.24 2.52 2.24
                 2.52 1.22 2.84 1.22 2.84 1.92 4.54 1.92 4.54 1.22 6.14 1.22
                 6.14 2.20 7.46 2.20 ;
        POLYGON  4.64 4.30 3.96 4.30 3.96 4.54 3.64 4.54 3.64 3.98 4.64 3.98 ;
        POLYGON  4.22 1.60 3.90 1.60 3.90 1.54 3.22 1.54 3.22 1.22 4.22 1.22 ;
        RECT  2.26 4.22 3.26 4.54 ;
        POLYGON  2.18 3.42 0.50 3.42 0.50 4.48 0.16 4.48 0.16 1.22 0.50 1.22
                 0.50 1.54 0.48 1.54 0.48 3.10 2.18 3.10 ;
    END
END latprs_4

MACRO latprs_2
    CLASS CORE ;
    FOREIGN latprs_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.76 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.72 3.68 3.36 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.58 2.72 14.26 2.72 14.26 2.40 14.24 2.40 14.24 2.08
                 14.58 2.08 ;
        END
    END gb
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.90  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  19.81 3.42 19.39 3.42 19.39 3.10 19.49 3.10 19.49 1.76
                 19.36 1.76 19.36 1.44 19.49 1.44 19.49 1.22 19.81 1.22 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.71  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  21.60 2.40 21.33 2.40 21.33 4.54 20.91 4.54 20.91 4.22
                 21.01 4.22 21.01 1.96 20.89 1.96 20.89 1.64 21.33 1.64
                 21.33 2.08 21.60 2.08 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  18.08 1.22 18.59 1.86 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.90  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.71 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.76 0.90 20.51 0.90 20.51 1.28 20.19 1.28 20.19 0.90
                 17.69 0.90 17.69 1.28 17.37 1.28 17.37 0.90 14.78 0.90
                 14.78 1.14 14.46 1.14 14.46 0.90 12.60 0.90 12.60 1.28
                 12.28 1.28 12.28 0.90 8.24 0.90 8.24 1.24 7.92 1.24 7.92 0.90
                 1.20 0.90 1.20 1.28 0.88 1.28 0.88 0.90 0.00 0.90 0.00 -0.90
                 21.76 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.76 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.16 1.20 4.16
                 1.20 4.86 1.56 4.86 1.56 4.16 1.88 4.16 1.88 4.86 12.28 4.86
                 12.28 4.16 12.60 4.16 12.60 4.86 14.42 4.86 14.42 4.16
                 15.30 4.16 15.30 4.86 16.67 4.86 16.67 2.95 16.99 2.95
                 16.99 4.86 21.76 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.67 2.62 20.59 2.62 20.59 4.54 17.43 4.54 17.43 2.52
                 16.21 2.52 16.21 3.21 15.89 3.21 15.89 2.18 15.46 2.18
                 15.28 2.00 15.28 1.22 15.60 1.22 15.60 1.86 16.21 1.86
                 16.21 2.20 17.75 2.20 17.75 4.22 20.27 4.22 20.27 2.30
                 20.67 2.30 ;
        RECT  18.71 2.76 19.05 3.90 ;
        RECT  15.98 1.22 16.99 1.54 ;
        POLYGON  15.22 3.84 5.34 3.84 5.34 4.30 5.02 4.30 5.02 3.52 5.18 3.52
                 5.18 1.90 5.50 1.90 5.50 3.52 14.90 3.52 14.90 2.40 15.22 2.40 ;
        POLYGON  14.08 1.54 13.94 1.54 13.94 1.95 13.82 2.07 13.82 2.48
                 13.94 2.60 13.94 2.88 13.98 2.88 13.98 3.20 13.62 3.20
                 13.62 2.74 13.50 2.62 13.50 1.93 13.62 1.81 13.62 1.22
                 14.08 1.22 ;
        POLYGON  13.30 1.62 13.18 1.74 13.18 2.88 13.30 2.88 13.30 3.20
                 6.16 3.20 6.16 2.88 12.86 2.88 12.86 1.47 12.91 1.47
                 12.91 1.37 12.98 1.37 12.98 1.30 13.30 1.30 ;
        POLYGON  11.92 1.60 11.60 1.60 11.60 1.54 8.88 1.54 8.88 1.88 7.28 1.88
                 7.28 1.60 6.46 1.60 6.46 1.28 7.60 1.28 7.60 1.56 8.56 1.56
                 8.56 1.22 11.92 1.22 ;
        POLYGON  11.92 4.54 5.72 4.54 5.72 4.16 6.04 4.16 6.04 4.22 11.92 4.22 ;
        POLYGON  11.22 2.52 8.70 2.52 8.70 2.20 10.90 2.20 10.90 2.04
                 11.22 2.04 ;
        POLYGON  7.46 2.52 5.82 2.52 5.82 1.54 4.86 1.54 4.86 2.24 2.52 2.24
                 2.52 1.22 2.84 1.22 2.84 1.92 4.54 1.92 4.54 1.22 6.14 1.22
                 6.14 2.20 7.46 2.20 ;
        POLYGON  4.64 4.30 3.96 4.30 3.96 4.54 3.64 4.54 3.64 3.98 4.64 3.98 ;
        POLYGON  4.22 1.60 3.90 1.60 3.90 1.54 3.22 1.54 3.22 1.22 4.22 1.22 ;
        RECT  2.26 4.22 3.26 4.54 ;
        POLYGON  2.18 3.42 0.50 3.42 0.50 4.48 0.16 4.48 0.16 1.22 0.50 1.22
                 0.50 1.54 0.48 1.54 0.48 3.10 2.18 3.10 ;
    END
END latprs_2

MACRO latprs_1
    CLASS CORE ;
    FOREIGN latprs_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.76 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.72 3.68 3.36 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.58 2.72 14.26 2.72 14.26 2.40 14.24 2.40 14.24 2.08
                 14.58 2.08 ;
        END
    END gb
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.46  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  19.81 3.66 19.39 3.66 19.39 3.34 19.49 3.34 19.49 1.76
                 19.36 1.76 19.36 1.44 19.49 1.44 19.49 1.22 19.81 1.22 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.23  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  21.60 2.40 21.33 2.40 21.33 4.54 20.91 4.54 20.91 4.22
                 21.01 4.22 21.01 1.54 20.89 1.54 20.89 1.22 21.33 1.22
                 21.33 2.08 21.60 2.08 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  18.08 1.22 18.59 1.86 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.90  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.71 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.76 0.90 20.51 0.90 20.51 1.26 20.19 1.26 20.19 0.90
                 17.69 0.90 17.69 1.28 17.37 1.28 17.37 0.90 14.78 0.90
                 14.78 1.14 14.46 1.14 14.46 0.90 12.60 0.90 12.60 1.28
                 12.28 1.28 12.28 0.90 8.24 0.90 8.24 1.24 7.92 1.24 7.92 0.90
                 1.20 0.90 1.20 1.28 0.88 1.28 0.88 0.90 0.00 0.90 0.00 -0.90
                 21.76 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.76 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.16 1.20 4.16
                 1.20 4.86 1.56 4.86 1.56 4.16 1.88 4.16 1.88 4.86 12.28 4.86
                 12.28 4.16 12.60 4.16 12.60 4.86 14.42 4.86 14.42 4.16
                 15.30 4.16 15.30 4.86 16.67 4.86 16.67 2.95 16.99 2.95
                 16.99 4.86 21.76 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.67 2.62 20.59 2.62 20.59 4.54 17.43 4.54 17.43 2.52
                 16.21 2.52 16.21 3.21 15.89 3.21 15.89 2.18 15.46 2.18
                 15.28 2.00 15.28 1.22 15.60 1.22 15.60 1.86 16.21 1.86
                 16.21 2.20 17.75 2.20 17.75 4.22 20.27 4.22 20.27 2.30
                 20.67 2.30 ;
        RECT  18.71 2.76 19.05 3.90 ;
        RECT  15.98 1.22 16.99 1.54 ;
        POLYGON  15.22 3.84 5.34 3.84 5.34 4.30 5.02 4.30 5.02 3.52 5.18 3.52
                 5.18 1.90 5.50 1.90 5.50 3.52 14.90 3.52 14.90 2.40 15.22 2.40 ;
        POLYGON  14.08 1.54 13.94 1.54 13.94 1.95 13.82 2.07 13.82 2.48
                 13.94 2.60 13.94 2.88 13.98 2.88 13.98 3.20 13.62 3.20
                 13.62 2.74 13.50 2.62 13.50 1.93 13.62 1.81 13.62 1.22
                 14.08 1.22 ;
        POLYGON  13.30 1.62 13.18 1.74 13.18 2.88 13.30 2.88 13.30 3.20
                 6.16 3.20 6.16 2.88 12.86 2.88 12.86 1.47 12.91 1.47
                 12.91 1.37 12.98 1.37 12.98 1.30 13.30 1.30 ;
        POLYGON  11.92 1.60 11.60 1.60 11.60 1.54 8.88 1.54 8.88 1.88 7.28 1.88
                 7.28 1.60 6.46 1.60 6.46 1.28 7.60 1.28 7.60 1.56 8.56 1.56
                 8.56 1.22 11.92 1.22 ;
        POLYGON  11.92 4.54 5.72 4.54 5.72 4.16 6.04 4.16 6.04 4.22 11.92 4.22 ;
        POLYGON  11.22 2.52 8.70 2.52 8.70 2.20 10.90 2.20 10.90 2.04
                 11.22 2.04 ;
        POLYGON  7.46 2.52 5.82 2.52 5.82 1.54 4.86 1.54 4.86 2.24 2.52 2.24
                 2.52 1.22 2.84 1.22 2.84 1.92 4.54 1.92 4.54 1.22 6.14 1.22
                 6.14 2.20 7.46 2.20 ;
        POLYGON  4.64 4.30 3.96 4.30 3.96 4.54 3.64 4.54 3.64 3.98 4.64 3.98 ;
        POLYGON  4.22 1.60 3.90 1.60 3.90 1.54 3.22 1.54 3.22 1.22 4.22 1.22 ;
        RECT  2.26 4.22 3.26 4.54 ;
        POLYGON  2.18 3.42 0.50 3.42 0.50 4.48 0.16 4.48 0.16 1.22 0.50 1.22
                 0.50 1.54 0.48 1.54 0.48 3.10 2.18 3.10 ;
    END
END latprs_1

MACRO latprqb_4
    CLASS CORE ;
    FOREIGN latprqb_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 13.44 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 4.00 2.57 4.46 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.82 3.04 ;
        END
    END gb
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  13.28 4.53 11.40 4.53 11.40 4.21 12.96 4.21 12.96 1.90
                 11.38 1.90 11.38 1.58 13.28 1.58 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.94 2.22 11.36 3.04 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  13.44 0.90 12.42 0.90 12.42 1.23 12.10 1.23 12.10 0.90
                 10.10 0.90 10.10 1.14 9.78 1.14 9.78 0.90 1.46 0.90 1.46 1.42
                 1.14 1.42 1.14 0.90 0.00 0.90 0.00 -0.90 13.44 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  13.44 6.66 0.00 6.66 0.00 4.86 1.14 4.86 1.14 4.14 1.46 4.14
                 1.46 4.86 13.44 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  12.42 3.89 11.04 3.89 11.04 3.95 10.72 3.95 10.72 3.89
                 8.98 3.89 8.98 3.26 8.46 3.26 8.46 2.94 9.30 2.94 9.30 3.57
                 10.30 3.57 10.30 1.40 10.48 1.22 10.80 1.22 10.80 1.54
                 10.62 1.54 10.62 3.57 12.10 3.57 12.10 2.34 12.42 2.34 ;
        POLYGON  9.94 3.00 9.62 3.00 9.62 2.52 8.14 2.52 8.14 3.58 8.66 3.58
                 8.66 4.22 9.40 4.22 9.40 4.54 8.34 4.54 8.34 3.90 6.68 3.90
                 6.54 4.04 6.54 4.54 6.22 4.54 6.22 3.90 6.54 3.58 7.82 3.58
                 7.82 2.52 7.08 2.52 6.32 1.76 6.32 1.22 6.64 1.22 6.64 1.62
                 7.22 2.20 9.94 2.20 ;
        RECT  8.40 1.22 9.40 1.54 ;
        RECT  7.02 1.22 8.02 1.54 ;
        RECT  6.92 4.22 8.02 4.54 ;
        POLYGON  6.06 3.24 5.40 3.90 4.30 3.90 4.30 4.54 3.28 4.54 3.28 4.22
                 3.98 4.22 3.98 3.58 5.26 3.58 5.74 3.10 5.74 2.50 5.42 2.18
                 2.70 2.18 2.70 1.86 5.56 1.86 6.06 2.36 ;
        RECT  4.94 1.22 5.94 1.54 ;
        RECT  4.84 4.22 5.84 4.54 ;
        POLYGON  5.42 2.96 3.66 2.96 3.66 3.68 0.76 3.68 0.76 3.86 0.44 3.86
                 0.44 3.36 1.14 3.36 1.14 2.18 0.36 2.18 0.36 1.86 1.46 1.86
                 1.46 3.36 3.34 3.36 3.34 2.64 5.42 2.64 ;
        POLYGON  4.56 1.54 2.38 1.54 2.38 2.58 2.92 2.58 2.92 2.90 2.06 2.90
                 2.06 1.22 4.56 1.22 ;
    END
END latprqb_4

MACRO latprqb_2
    CLASS CORE ;
    FOREIGN latprqb_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.80 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 4.00 2.57 4.46 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.82 3.04 ;
        END
    END gb
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.64 4.54 12.30 4.54 12.30 4.22 12.32 4.22 12.32 1.54
                 12.30 1.54 12.30 1.22 12.64 1.22 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  11.04 1.94 11.36 2.58 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  12.80 0.90 10.10 0.90 10.10 1.14 9.78 1.14 9.78 0.90 1.46 0.90
                 1.46 1.42 1.14 1.42 1.14 0.90 0.00 0.90 0.00 -0.90 12.80 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  12.80 6.66 0.00 6.66 0.00 4.86 1.14 4.86 1.14 4.14 1.46 4.14
                 1.46 4.86 12.80 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  12.00 3.74 11.20 4.54 10.40 4.54 10.40 3.90 8.98 3.90
                 8.98 3.26 8.46 3.26 8.46 2.94 9.30 2.94 9.30 3.58 10.40 3.58
                 10.40 1.30 10.48 1.22 10.80 1.22 10.80 1.54 10.72 1.54
                 10.72 4.22 11.05 4.22 11.68 3.59 11.68 2.14 12.00 2.14 ;
        POLYGON  9.94 3.00 9.62 3.00 9.62 2.52 8.14 2.52 8.14 3.58 8.66 3.58
                 8.66 4.22 9.40 4.22 9.40 4.54 8.34 4.54 8.34 3.90 6.68 3.90
                 6.54 4.04 6.54 4.54 6.22 4.54 6.22 3.90 6.54 3.58 7.82 3.58
                 7.82 2.52 7.08 2.52 6.32 1.76 6.32 1.22 6.64 1.22 6.64 1.62
                 7.22 2.20 9.94 2.20 ;
        RECT  8.40 1.22 9.40 1.54 ;
        RECT  7.02 1.22 8.02 1.54 ;
        RECT  6.92 4.22 8.02 4.54 ;
        POLYGON  6.06 3.24 5.40 3.90 4.30 3.90 4.30 4.54 3.28 4.54 3.28 4.22
                 3.98 4.22 3.98 3.58 5.26 3.58 5.74 3.10 5.74 2.50 5.42 2.18
                 2.70 2.18 2.70 1.86 5.56 1.86 6.06 2.36 ;
        RECT  4.94 1.22 5.94 1.54 ;
        RECT  4.84 4.22 5.84 4.54 ;
        POLYGON  5.42 2.96 3.66 2.96 3.66 3.68 0.76 3.68 0.76 3.86 0.44 3.86
                 0.44 3.36 1.14 3.36 1.14 2.18 0.36 2.18 0.36 1.86 1.46 1.86
                 1.46 3.36 3.34 3.36 3.34 2.64 5.42 2.64 ;
        POLYGON  4.56 1.54 2.38 1.54 2.38 2.58 2.92 2.58 2.92 2.90 2.06 2.90
                 2.06 1.22 4.56 1.22 ;
    END
END latprqb_2

MACRO latprqb_1
    CLASS CORE ;
    FOREIGN latprqb_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.80 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 4.00 2.57 4.46 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.82 3.04 ;
        END
    END gb
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.64 4.54 12.30 4.54 12.30 4.22 12.32 4.22 12.32 1.54
                 12.30 1.54 12.30 1.22 12.64 1.22 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  11.04 1.94 11.36 2.58 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  12.80 0.90 10.10 0.90 10.10 1.14 9.78 1.14 9.78 0.90 1.46 0.90
                 1.46 1.42 1.14 1.42 1.14 0.90 0.00 0.90 0.00 -0.90 12.80 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  12.80 6.66 0.00 6.66 0.00 4.86 1.14 4.86 1.14 4.14 1.46 4.14
                 1.46 4.86 12.80 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  12.00 3.74 11.20 4.54 10.40 4.54 10.40 3.90 8.98 3.90
                 8.98 3.26 8.46 3.26 8.46 2.94 9.30 2.94 9.30 3.58 10.40 3.58
                 10.40 1.30 10.48 1.22 10.80 1.22 10.80 1.54 10.72 1.54
                 10.72 4.22 11.05 4.22 11.68 3.59 11.68 2.14 12.00 2.14 ;
        POLYGON  9.94 3.00 9.62 3.00 9.62 2.52 8.14 2.52 8.14 3.58 8.66 3.58
                 8.66 4.22 9.40 4.22 9.40 4.54 8.34 4.54 8.34 3.90 6.68 3.90
                 6.54 4.04 6.54 4.54 6.22 4.54 6.22 3.90 6.54 3.58 7.82 3.58
                 7.82 2.52 7.08 2.52 6.32 1.76 6.32 1.22 6.64 1.22 6.64 1.62
                 7.22 2.20 9.94 2.20 ;
        RECT  8.40 1.22 9.40 1.54 ;
        RECT  7.02 1.22 8.02 1.54 ;
        RECT  6.92 4.22 8.02 4.54 ;
        POLYGON  6.06 3.24 5.40 3.90 4.30 3.90 4.30 4.54 3.28 4.54 3.28 4.22
                 3.98 4.22 3.98 3.58 5.26 3.58 5.74 3.10 5.74 2.50 5.42 2.18
                 2.70 2.18 2.70 1.86 5.56 1.86 6.06 2.36 ;
        RECT  4.94 1.22 5.94 1.54 ;
        RECT  4.84 4.22 5.84 4.54 ;
        POLYGON  5.42 2.96 3.66 2.96 3.66 3.68 0.76 3.68 0.76 3.86 0.44 3.86
                 0.44 3.36 1.14 3.36 1.14 2.18 0.36 2.18 0.36 1.86 1.46 1.86
                 1.46 3.36 3.34 3.36 3.34 2.64 5.42 2.64 ;
        POLYGON  4.56 1.54 2.38 1.54 2.38 2.58 2.92 2.58 2.92 2.90 2.06 2.90
                 2.06 1.22 4.56 1.22 ;
    END
END latprqb_1

MACRO latprq_4
    CLASS CORE ;
    FOREIGN latprq_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.08 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 4.00 2.57 4.46 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.82 3.04 ;
        END
    END gb
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  13.63 3.25 11.86 3.25 11.86 2.93 12.96 2.93 12.96 2.71
                 13.31 2.71 13.31 1.62 11.38 1.62 11.38 1.30 13.63 1.30 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.94 1.94 11.36 2.58 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  14.08 0.90 10.10 0.90 10.10 1.14 9.78 1.14 9.78 0.90 1.46 0.90
                 1.46 1.42 1.14 1.42 1.14 0.90 0.00 0.90 0.00 -0.90 14.08 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  14.08 6.66 0.00 6.66 0.00 4.86 1.14 4.86 1.14 4.14 1.46 4.14
                 1.46 4.86 12.50 4.86 12.50 4.79 12.92 4.79 12.92 4.86
                 14.08 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  11.04 4.37 10.30 4.37 10.30 3.90 8.98 3.90 8.98 3.26 8.46 3.26
                 8.46 2.94 9.30 2.94 9.30 3.58 10.30 3.58 10.30 1.40 10.48 1.22
                 10.80 1.22 10.80 1.54 10.62 1.54 10.62 4.05 11.04 4.05 ;
        POLYGON  9.94 3.00 9.62 3.00 9.62 2.52 8.14 2.52 8.14 3.58 8.66 3.58
                 8.66 4.22 9.40 4.22 9.40 4.54 8.34 4.54 8.34 3.90 6.68 3.90
                 6.54 4.04 6.54 4.54 6.22 4.54 6.22 3.90 6.54 3.58 7.82 3.58
                 7.82 2.52 7.08 2.52 6.32 1.76 6.32 1.22 6.64 1.22 6.64 1.62
                 7.22 2.20 9.94 2.20 ;
        RECT  8.40 1.22 9.40 1.54 ;
        RECT  7.02 1.22 8.02 1.54 ;
        RECT  6.92 4.22 8.02 4.54 ;
        POLYGON  6.06 3.24 5.40 3.90 4.30 3.90 4.30 4.54 3.28 4.54 3.28 4.22
                 3.98 4.22 3.98 3.58 5.26 3.58 5.74 3.10 5.74 2.50 5.42 2.18
                 2.70 2.18 2.70 1.86 5.56 1.86 6.06 2.36 ;
        RECT  4.94 1.22 5.94 1.54 ;
        RECT  4.84 4.22 5.84 4.54 ;
        POLYGON  5.42 2.96 3.66 2.96 3.66 3.68 0.76 3.68 0.76 3.86 0.44 3.86
                 0.44 3.36 1.14 3.36 1.14 2.18 0.36 2.18 0.36 1.86 1.46 1.86
                 1.46 3.36 3.34 3.36 3.34 2.64 5.42 2.64 ;
        POLYGON  4.56 1.54 2.38 1.54 2.38 2.58 2.92 2.58 2.92 2.90 2.06 2.90
                 2.06 1.22 4.56 1.22 ;
    END
END latprq_4

MACRO latprq_2
    CLASS CORE ;
    FOREIGN latprq_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.80 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 4.00 2.57 4.46 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.82 3.04 ;
        END
    END gb
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.64 3.04 12.42 3.04 12.42 4.54 12.10 4.54 12.10 1.64
                 12.42 1.64 12.42 2.72 12.64 2.72 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  11.04 2.08 11.36 2.89 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  12.80 0.90 11.72 0.90 11.72 1.42 11.40 1.42 11.40 0.90
                 10.10 0.90 10.10 1.14 9.78 1.14 9.78 0.90 1.46 0.90 1.46 1.42
                 1.14 1.42 1.14 0.90 0.00 0.90 0.00 -0.90 12.80 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  12.80 6.66 0.00 6.66 0.00 4.86 1.14 4.86 1.14 4.14 1.46 4.14
                 1.46 4.86 11.40 4.86 11.40 4.22 11.72 4.22 11.72 4.86
                 12.80 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  11.04 4.54 10.40 4.54 10.40 3.90 8.98 3.90 8.98 3.26 8.46 3.26
                 8.46 2.94 9.30 2.94 9.30 3.58 10.40 3.58 10.40 1.30 10.48 1.22
                 10.80 1.22 10.80 1.54 10.72 1.54 10.72 4.22 11.04 4.22 ;
        POLYGON  9.94 3.00 9.62 3.00 9.62 2.52 8.14 2.52 8.14 3.58 8.66 3.58
                 8.66 4.22 9.40 4.22 9.40 4.54 8.34 4.54 8.34 3.90 6.68 3.90
                 6.54 4.04 6.54 4.54 6.22 4.54 6.22 3.90 6.54 3.58 7.82 3.58
                 7.82 2.52 7.08 2.52 6.32 1.76 6.32 1.22 6.64 1.22 6.64 1.62
                 7.22 2.20 9.94 2.20 ;
        RECT  8.40 1.22 9.40 1.54 ;
        RECT  7.02 1.22 8.02 1.54 ;
        RECT  6.92 4.22 8.02 4.54 ;
        POLYGON  6.06 3.24 5.40 3.90 4.30 3.90 4.30 4.54 3.28 4.54 3.28 4.22
                 3.98 4.22 3.98 3.58 5.26 3.58 5.74 3.10 5.74 2.50 5.42 2.18
                 2.70 2.18 2.70 1.86 5.56 1.86 6.06 2.36 ;
        RECT  4.94 1.22 5.94 1.54 ;
        RECT  4.84 4.22 5.84 4.54 ;
        POLYGON  5.42 2.96 3.66 2.96 3.66 3.68 0.76 3.68 0.76 3.86 0.44 3.86
                 0.44 3.36 1.14 3.36 1.14 2.18 0.36 2.18 0.36 1.86 1.46 1.86
                 1.46 3.36 3.34 3.36 3.34 2.64 5.42 2.64 ;
        POLYGON  4.56 1.54 2.38 1.54 2.38 2.58 2.92 2.58 2.92 2.90 2.06 2.90
                 2.06 1.22 4.56 1.22 ;
    END
END latprq_2

MACRO latprq_1
    CLASS CORE ;
    FOREIGN latprq_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.80 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 4.00 2.57 4.46 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.82 3.04 ;
        END
    END gb
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.64 3.04 12.42 3.04 12.42 4.54 12.10 4.54 12.10 1.22
                 12.42 1.22 12.42 2.72 12.64 2.72 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  11.04 1.94 11.36 2.58 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  12.80 0.90 11.72 0.90 11.72 1.54 11.40 1.54 11.40 0.90
                 10.10 0.90 10.10 1.14 9.78 1.14 9.78 0.90 1.46 0.90 1.46 1.42
                 1.14 1.42 1.14 0.90 0.00 0.90 0.00 -0.90 12.80 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  12.80 6.66 0.00 6.66 0.00 4.86 1.14 4.86 1.14 4.14 1.46 4.14
                 1.46 4.86 11.40 4.86 11.40 4.22 11.72 4.22 11.72 4.86
                 12.80 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  11.04 4.54 10.40 4.54 10.40 3.90 8.98 3.90 8.98 3.26 8.46 3.26
                 8.46 2.94 9.30 2.94 9.30 3.58 10.40 3.58 10.40 1.30 10.48 1.22
                 10.80 1.22 10.80 1.54 10.72 1.54 10.72 4.22 11.04 4.22 ;
        POLYGON  9.94 3.00 9.62 3.00 9.62 2.52 8.14 2.52 8.14 3.58 8.66 3.58
                 8.66 4.22 9.40 4.22 9.40 4.54 8.34 4.54 8.34 3.90 6.68 3.90
                 6.54 4.04 6.54 4.54 6.22 4.54 6.22 3.90 6.54 3.58 7.82 3.58
                 7.82 2.52 7.08 2.52 6.32 1.76 6.32 1.22 6.64 1.22 6.64 1.62
                 7.22 2.20 9.94 2.20 ;
        RECT  8.40 1.22 9.40 1.54 ;
        RECT  7.02 1.22 8.02 1.54 ;
        RECT  6.92 4.22 8.02 4.54 ;
        POLYGON  6.06 3.24 5.40 3.90 4.30 3.90 4.30 4.54 3.28 4.54 3.28 4.22
                 3.98 4.22 3.98 3.58 5.26 3.58 5.74 3.10 5.74 2.50 5.42 2.18
                 2.70 2.18 2.70 1.86 5.56 1.86 6.06 2.36 ;
        RECT  4.94 1.22 5.94 1.54 ;
        RECT  4.84 4.22 5.84 4.54 ;
        POLYGON  5.42 2.96 3.66 2.96 3.66 3.68 0.76 3.68 0.76 3.86 0.44 3.86
                 0.44 3.36 1.14 3.36 1.14 2.18 0.36 2.18 0.36 1.86 1.46 1.86
                 1.46 3.36 3.34 3.36 3.34 2.64 5.42 2.64 ;
        POLYGON  4.56 1.54 2.38 1.54 2.38 2.58 2.92 2.58 2.92 2.90 2.06 2.90
                 2.06 1.22 4.56 1.22 ;
    END
END latprq_1

MACRO latpr_4
    CLASS CORE ;
    FOREIGN latpr_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.00 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 4.00 2.57 4.46 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.82 3.04 ;
        END
    END gb
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  13.63 3.25 11.86 3.25 11.86 2.93 12.96 2.93 12.96 2.72
                 13.31 2.72 13.31 1.62 11.38 1.62 11.38 1.30 13.63 1.30 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  15.84 4.53 13.95 4.53 13.95 4.21 15.52 4.21 15.52 1.90
                 13.95 1.90 13.95 1.58 15.84 1.58 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.94 1.94 11.36 2.58 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 0.90 14.97 0.90 14.97 1.23 14.65 1.23 14.65 0.90
                 10.10 0.90 10.10 1.14 9.78 1.14 9.78 0.90 1.46 0.90 1.46 1.42
                 1.14 1.42 1.14 0.90 0.00 0.90 0.00 -0.90 16.00 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 6.66 0.00 6.66 0.00 4.86 1.14 4.86 1.14 4.14 1.46 4.14
                 1.46 4.86 12.50 4.86 12.50 4.79 12.92 4.79 12.92 4.86
                 16.00 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  14.97 3.89 12.64 3.89 12.64 4.37 10.30 4.37 10.30 3.90
                 8.98 3.90 8.98 3.26 8.46 3.26 8.46 2.94 9.30 2.94 9.30 3.58
                 10.30 3.58 10.30 1.40 10.48 1.22 10.80 1.22 10.80 1.54
                 10.62 1.54 10.62 4.05 12.32 4.05 12.32 3.57 14.65 3.57
                 14.65 2.34 14.97 2.34 ;
        POLYGON  9.94 3.00 9.62 3.00 9.62 2.52 8.14 2.52 8.14 3.58 8.66 3.58
                 8.66 4.22 9.40 4.22 9.40 4.54 8.34 4.54 8.34 3.90 6.68 3.90
                 6.54 4.04 6.54 4.54 6.22 4.54 6.22 3.90 6.54 3.58 7.82 3.58
                 7.82 2.52 7.08 2.52 6.32 1.76 6.32 1.22 6.64 1.22 6.64 1.62
                 7.22 2.20 9.94 2.20 ;
        RECT  8.40 1.22 9.40 1.54 ;
        RECT  7.02 1.22 8.02 1.54 ;
        RECT  6.92 4.22 8.02 4.54 ;
        POLYGON  6.06 3.24 5.40 3.90 4.30 3.90 4.30 4.54 3.28 4.54 3.28 4.22
                 3.98 4.22 3.98 3.58 5.26 3.58 5.74 3.10 5.74 2.50 5.42 2.18
                 2.70 2.18 2.70 1.86 5.56 1.86 6.06 2.36 ;
        RECT  4.94 1.22 5.94 1.54 ;
        RECT  4.84 4.22 5.84 4.54 ;
        POLYGON  5.42 2.96 3.66 2.96 3.66 3.68 0.76 3.68 0.76 3.86 0.44 3.86
                 0.44 3.36 1.14 3.36 1.14 2.18 0.36 2.18 0.36 1.86 1.46 1.86
                 1.46 3.36 3.34 3.36 3.34 2.64 5.42 2.64 ;
        POLYGON  4.56 1.54 2.38 1.54 2.38 2.58 2.92 2.58 2.92 2.90 2.06 2.90
                 2.06 1.22 4.56 1.22 ;
    END
END latpr_4

MACRO latpr_2
    CLASS CORE ;
    FOREIGN latpr_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 13.44 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 4.00 2.57 4.46 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.82 3.04 ;
        END
    END gb
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.99  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.00 3.40 11.40 3.40 11.40 3.08 11.58 3.08 11.68 2.98
                 11.68 1.57 11.40 1.57 11.40 1.25 12.00 1.25 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  13.28 4.54 12.94 4.54 12.94 4.22 12.96 4.22 12.96 1.96
                 12.94 1.96 12.94 1.64 13.28 1.64 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  11.04 2.08 11.36 2.73 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  13.44 0.90 10.10 0.90 10.10 1.14 9.78 1.14 9.78 0.90 1.46 0.90
                 1.46 1.42 1.14 1.42 1.14 0.90 0.00 0.90 0.00 -0.90 13.44 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  13.44 6.66 0.00 6.66 0.00 4.86 1.14 4.86 1.14 4.14 1.46 4.14
                 1.46 4.86 13.44 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  12.64 3.90 12.00 4.54 10.40 4.54 10.40 3.90 8.98 3.90
                 8.98 3.26 8.46 3.26 8.46 2.94 9.30 2.94 9.30 3.58 10.40 3.58
                 10.40 1.30 10.48 1.22 10.80 1.22 10.80 1.54 10.72 1.54
                 10.72 4.22 11.86 4.22 12.32 3.76 12.32 2.14 12.64 2.14 ;
        POLYGON  9.94 3.00 9.62 3.00 9.62 2.52 8.14 2.52 8.14 3.58 8.66 3.58
                 8.66 4.22 9.40 4.22 9.40 4.54 8.34 4.54 8.34 3.90 6.68 3.90
                 6.54 4.04 6.54 4.54 6.22 4.54 6.22 3.90 6.54 3.58 7.82 3.58
                 7.82 2.52 7.08 2.52 6.32 1.76 6.32 1.22 6.64 1.22 6.64 1.62
                 7.22 2.20 9.94 2.20 ;
        RECT  8.40 1.22 9.40 1.54 ;
        RECT  7.02 1.22 8.02 1.54 ;
        RECT  6.92 4.22 8.02 4.54 ;
        POLYGON  6.06 3.24 5.40 3.90 4.30 3.90 4.30 4.54 3.28 4.54 3.28 4.22
                 3.98 4.22 3.98 3.58 5.26 3.58 5.74 3.10 5.74 2.50 5.42 2.18
                 2.70 2.18 2.70 1.86 5.56 1.86 6.06 2.36 ;
        RECT  4.94 1.22 5.94 1.54 ;
        RECT  4.84 4.22 5.84 4.54 ;
        POLYGON  5.42 2.96 3.66 2.96 3.66 3.68 0.76 3.68 0.76 3.86 0.44 3.86
                 0.44 3.36 1.14 3.36 1.14 2.18 0.36 2.18 0.36 1.86 1.46 1.86
                 1.46 3.36 3.34 3.36 3.34 2.64 5.42 2.64 ;
        POLYGON  4.56 1.54 2.38 1.54 2.38 2.58 2.92 2.58 2.92 2.90 2.06 2.90
                 2.06 1.22 4.56 1.22 ;
    END
END latpr_2

MACRO latpr_1
    CLASS CORE ;
    FOREIGN latpr_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 13.44 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 4.00 2.57 4.46 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.82 3.04 ;
        END
    END gb
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.00 3.38 11.72 3.66 11.40 3.66 11.40 3.34 11.58 3.34
                 11.68 3.24 11.68 1.54 11.40 1.54 11.40 1.22 12.00 1.22 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  13.28 4.54 12.94 4.54 12.94 4.22 12.96 4.22 12.96 1.54
                 12.94 1.54 12.94 1.22 13.28 1.22 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  11.04 1.94 11.36 2.58 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  13.44 0.90 10.10 0.90 10.10 1.14 9.78 1.14 9.78 0.90 1.46 0.90
                 1.46 1.42 1.14 1.42 1.14 0.90 0.00 0.90 0.00 -0.90 13.44 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  13.44 6.66 0.00 6.66 0.00 4.86 1.14 4.86 1.14 4.14 1.46 4.14
                 1.46 4.86 13.44 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  12.64 3.90 12.00 4.54 10.40 4.54 10.40 3.90 8.98 3.90
                 8.98 3.26 8.46 3.26 8.46 2.94 9.30 2.94 9.30 3.58 10.40 3.58
                 10.40 1.30 10.48 1.22 10.80 1.22 10.80 1.54 10.72 1.54
                 10.72 4.22 11.86 4.22 12.32 3.76 12.32 2.14 12.64 2.14 ;
        POLYGON  9.94 3.00 9.62 3.00 9.62 2.52 8.14 2.52 8.14 3.58 8.66 3.58
                 8.66 4.22 9.40 4.22 9.40 4.54 8.34 4.54 8.34 3.90 6.68 3.90
                 6.54 4.04 6.54 4.54 6.22 4.54 6.22 3.90 6.54 3.58 7.82 3.58
                 7.82 2.52 7.08 2.52 6.32 1.76 6.32 1.22 6.64 1.22 6.64 1.62
                 7.22 2.20 9.94 2.20 ;
        RECT  8.40 1.22 9.40 1.54 ;
        RECT  7.02 1.22 8.02 1.54 ;
        RECT  6.92 4.22 8.02 4.54 ;
        POLYGON  6.06 3.24 5.40 3.90 4.30 3.90 4.30 4.54 3.28 4.54 3.28 4.22
                 3.98 4.22 3.98 3.58 5.26 3.58 5.74 3.10 5.74 2.50 5.42 2.18
                 2.70 2.18 2.70 1.86 5.56 1.86 6.06 2.36 ;
        RECT  4.94 1.22 5.94 1.54 ;
        RECT  4.84 4.22 5.84 4.54 ;
        POLYGON  5.42 2.96 3.66 2.96 3.66 3.68 0.76 3.68 0.76 3.86 0.44 3.86
                 0.44 3.36 1.14 3.36 1.14 2.18 0.36 2.18 0.36 1.86 1.46 1.86
                 1.46 3.36 3.34 3.36 3.34 2.64 5.42 2.64 ;
        POLYGON  4.56 1.54 2.38 1.54 2.38 2.58 2.92 2.58 2.92 2.90 2.06 2.90
                 2.06 1.22 4.56 1.22 ;
    END
END latpr_1

MACRO latpqb_4
    CLASS CORE ;
    FOREIGN latpqb_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.88 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.16 4.53 8.44 4.53 8.44 4.21 9.84 4.21 9.84 3.04 9.76 3.04
                 9.76 2.72 9.84 2.72 9.84 1.90 8.44 1.90 8.44 1.58 10.16 1.58 ;
        END
    END qb
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.08 7.12 2.54 ;
        END
    END gb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  10.88 0.90 9.46 0.90 9.46 1.23 9.14 1.23 9.14 0.90 7.06 0.90
                 7.06 1.12 6.74 1.12 6.74 0.90 4.88 0.90 4.88 1.14 4.56 1.14
                 4.56 0.90 1.20 0.90 1.20 1.62 0.88 1.62 0.88 0.90 0.00 0.90
                 0.00 -0.90 10.88 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  10.88 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 4.66 4.86 4.66 4.62 4.98 4.62 4.98 4.86 6.74 4.86
                 6.74 4.62 7.06 4.62 7.06 4.86 10.88 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  9.44 3.58 8.12 3.58 8.12 4.54 7.80 4.54 7.80 3.74 7.44 3.74
                 7.44 3.42 7.54 3.42 7.54 2.11 7.44 2.11 7.44 1.22 7.76 1.22
                 7.76 1.83 7.86 1.83 7.86 3.26 9.12 3.26 9.12 2.34 9.44 2.34 ;
        POLYGON  7.22 3.18 7.00 3.18 7.00 4.30 4.66 4.30 4.66 3.90 2.80 3.90
                 2.80 4.54 2.48 4.54 2.48 1.30 2.80 1.30 2.80 3.58 4.98 3.58
                 4.98 3.98 6.68 3.98 6.68 2.86 7.22 2.86 ;
        POLYGON  6.36 1.54 6.32 1.54 6.32 1.80 5.97 2.15 5.97 2.71 6.32 3.06
                 6.32 3.34 6.36 3.34 6.36 3.66 6.00 3.66 6.00 3.20 5.65 2.85
                 5.65 2.01 6.00 1.66 6.00 1.22 6.36 1.22 ;
        POLYGON  5.68 3.66 5.36 3.66 5.36 3.48 5.14 3.26 4.66 3.26 4.66 2.58
                 3.70 2.58 3.70 2.26 4.66 2.26 4.66 1.90 5.26 1.30 5.58 1.30
                 5.58 1.62 5.40 1.62 4.98 2.04 4.98 2.94 5.28 2.94 5.68 3.34 ;
        RECT  3.18 4.22 4.28 4.54 ;
        RECT  3.18 1.58 4.18 1.90 ;
        POLYGON  2.00 2.26 0.18 2.26 0.18 1.30 0.50 1.30 0.50 1.94 1.68 1.94
                 1.68 1.30 2.00 1.30 ;
        POLYGON  1.88 4.54 1.56 4.54 1.56 3.76 0.50 3.76 0.50 4.54 0.18 4.54
                 0.18 3.44 1.88 3.44 ;
    END
END latpqb_4

MACRO latpqb_2
    CLASS CORE ;
    FOREIGN latpqb_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.60 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.08 7.16 2.54 ;
        END
    END gb
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.44 4.30 8.94 4.30 8.94 3.98 9.12 3.98 9.12 1.96 8.94 1.96
                 8.94 1.64 9.44 1.64 ;
        END
    END qb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  9.60 0.90 8.56 0.90 8.56 1.08 8.24 1.08 8.24 0.90 7.06 0.90
                 7.06 1.12 6.74 1.12 6.74 0.90 4.88 0.90 4.88 1.14 4.56 1.14
                 4.56 0.90 1.20 0.90 1.20 1.62 0.88 1.62 0.88 0.90 0.00 0.90
                 0.00 -0.90 9.60 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  9.60 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 4.66 4.86 4.66 4.62 4.98 4.62 4.98 4.86 6.74 4.86
                 6.74 4.62 7.06 4.62 7.06 4.86 9.60 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  8.72 2.62 7.86 2.62 7.86 3.78 8.12 3.78 8.12 4.54 7.80 4.54
                 7.80 4.10 7.54 4.10 7.54 3.74 7.44 3.74 7.44 3.42 7.54 3.42
                 7.54 1.54 7.44 1.54 7.44 1.22 7.86 1.22 7.86 2.30 8.72 2.30 ;
        POLYGON  7.22 3.18 7.00 3.18 7.00 4.30 4.66 4.30 4.66 3.90 2.80 3.90
                 2.80 4.54 2.48 4.54 2.48 1.30 2.80 1.30 2.80 3.58 4.98 3.58
                 4.98 3.98 6.68 3.98 6.68 2.86 7.22 2.86 ;
        POLYGON  6.36 1.54 6.32 1.54 6.32 1.80 5.97 2.15 5.97 2.71 6.32 3.06
                 6.32 3.34 6.36 3.34 6.36 3.66 6.00 3.66 6.00 3.20 5.65 2.85
                 5.65 2.01 6.00 1.66 6.00 1.22 6.36 1.22 ;
        POLYGON  5.68 3.66 5.36 3.66 5.36 3.48 5.14 3.26 4.66 3.26 4.66 2.58
                 3.70 2.58 3.70 2.26 4.66 2.26 4.66 1.90 5.26 1.30 5.58 1.30
                 5.58 1.62 5.40 1.62 4.98 2.04 4.98 2.94 5.28 2.94 5.68 3.34 ;
        RECT  3.18 4.22 4.28 4.54 ;
        RECT  3.18 1.58 4.18 1.90 ;
        POLYGON  2.00 2.26 0.18 2.26 0.18 1.30 0.50 1.30 0.50 1.94 1.68 1.94
                 1.68 1.30 2.00 1.30 ;
        POLYGON  1.88 4.54 1.56 4.54 1.56 3.76 0.50 3.76 0.50 4.54 0.18 4.54
                 0.18 3.44 1.88 3.44 ;
    END
END latpqb_2

MACRO latpqb_1
    CLASS CORE ;
    FOREIGN latpqb_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.60 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.08 7.16 2.54 ;
        END
    END gb
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.44 4.30 8.94 4.30 8.94 3.98 9.12 3.98 9.12 1.54 8.94 1.54
                 8.94 1.22 9.44 1.22 ;
        END
    END qb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  9.60 0.90 8.56 0.90 8.56 1.08 8.24 1.08 8.24 0.90 7.06 0.90
                 7.06 1.12 6.74 1.12 6.74 0.90 4.88 0.90 4.88 1.14 4.56 1.14
                 4.56 0.90 1.20 0.90 1.20 1.62 0.88 1.62 0.88 0.90 0.00 0.90
                 0.00 -0.90 9.60 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  9.60 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 4.66 4.86 4.66 4.62 4.98 4.62 4.98 4.86 6.74 4.86
                 6.74 4.62 7.06 4.62 7.06 4.86 9.60 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  8.72 2.62 7.86 2.62 7.86 3.78 8.12 3.78 8.12 4.54 7.80 4.54
                 7.80 4.10 7.54 4.10 7.54 3.74 7.44 3.74 7.44 3.42 7.54 3.42
                 7.54 1.54 7.44 1.54 7.44 1.22 7.86 1.22 7.86 2.30 8.72 2.30 ;
        POLYGON  7.22 3.18 7.00 3.18 7.00 4.30 4.66 4.30 4.66 3.90 2.80 3.90
                 2.80 4.54 2.48 4.54 2.48 1.30 2.80 1.30 2.80 3.58 4.98 3.58
                 4.98 3.98 6.68 3.98 6.68 2.86 7.22 2.86 ;
        POLYGON  6.36 1.54 6.32 1.54 6.32 1.80 5.97 2.15 5.97 2.71 6.32 3.06
                 6.32 3.34 6.36 3.34 6.36 3.66 6.00 3.66 6.00 3.20 5.65 2.85
                 5.65 2.01 6.00 1.66 6.00 1.22 6.36 1.22 ;
        POLYGON  5.68 3.66 5.36 3.66 5.36 3.48 5.14 3.26 4.66 3.26 4.66 2.58
                 3.70 2.58 3.70 2.26 4.66 2.26 4.66 1.90 5.26 1.30 5.58 1.30
                 5.58 1.62 5.40 1.62 4.98 2.04 4.98 2.94 5.28 2.94 5.68 3.34 ;
        RECT  3.18 4.22 4.28 4.54 ;
        RECT  3.18 1.58 4.18 1.90 ;
        POLYGON  2.00 2.26 0.18 2.26 0.18 1.30 0.50 1.30 0.50 1.94 1.68 1.94
                 1.68 1.30 2.00 1.30 ;
        POLYGON  1.88 4.54 1.56 4.54 1.56 3.76 0.50 3.76 0.50 4.54 0.18 4.54
                 0.18 3.44 1.88 3.44 ;
    END
END latpqb_1

MACRO latpq_4
    CLASS CORE ;
    FOREIGN latpq_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.88 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.08 7.12 2.54 ;
        END
    END gb
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.37 3.25 8.60 3.25 8.60 2.93 9.76 2.93 9.76 2.72 10.05 2.72
                 10.05 1.62 8.12 1.62 8.12 1.30 10.37 1.30 ;
        END
    END q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  10.88 0.90 7.06 0.90 7.06 1.12 6.74 1.12 6.74 0.90 4.88 0.90
                 4.88 1.14 4.56 1.14 4.56 0.90 1.20 0.90 1.20 1.62 0.88 1.62
                 0.88 0.90 0.00 0.90 0.00 -0.90 10.88 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  10.88 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 4.66 4.86 4.66 4.62 4.98 4.62 4.98 4.86 6.74 4.86
                 6.74 4.62 7.06 4.62 7.06 4.86 9.24 4.86 9.24 4.79 9.66 4.79
                 9.66 4.86 10.88 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  8.12 4.54 7.80 4.54 7.80 4.10 7.54 4.10 7.54 3.74 7.44 3.74
                 7.44 3.42 7.54 3.42 7.54 2.11 7.44 2.11 7.44 1.22 7.76 1.22
                 7.76 1.83 7.86 1.83 7.86 3.78 8.12 3.78 ;
        POLYGON  7.22 3.18 7.00 3.18 7.00 4.30 4.66 4.30 4.66 3.90 2.80 3.90
                 2.80 4.54 2.48 4.54 2.48 1.30 2.80 1.30 2.80 3.58 4.98 3.58
                 4.98 3.98 6.68 3.98 6.68 2.86 7.22 2.86 ;
        POLYGON  6.36 1.54 6.32 1.54 6.32 1.80 5.97 2.15 5.97 2.71 6.32 3.06
                 6.32 3.34 6.36 3.34 6.36 3.66 6.00 3.66 6.00 3.20 5.65 2.85
                 5.65 2.01 6.00 1.66 6.00 1.22 6.36 1.22 ;
        POLYGON  5.68 3.66 5.36 3.66 5.36 3.48 5.14 3.26 4.66 3.26 4.66 2.58
                 3.70 2.58 3.70 2.26 4.66 2.26 4.66 1.90 5.26 1.30 5.58 1.30
                 5.58 1.62 5.40 1.62 4.98 2.04 4.98 2.94 5.28 2.94 5.68 3.34 ;
        RECT  3.18 4.22 4.28 4.54 ;
        RECT  3.18 1.58 4.18 1.90 ;
        POLYGON  2.00 2.26 0.18 2.26 0.18 1.30 0.50 1.30 0.50 1.94 1.68 1.94
                 1.68 1.30 2.00 1.30 ;
        POLYGON  1.88 4.54 1.56 4.54 1.56 3.76 0.50 3.76 0.50 4.54 0.18 4.54
                 0.18 3.44 1.88 3.44 ;
    END
END latpq_4

MACRO latpq_2
    CLASS CORE ;
    FOREIGN latpq_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.60 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.08 7.16 2.54 ;
        END
    END gb
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.44 2.40 9.26 2.40 9.26 4.54 8.94 4.54 8.94 1.64 9.26 1.64
                 9.26 2.08 9.44 2.08 ;
        END
    END q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  9.60 0.90 8.56 0.90 8.56 1.96 8.24 1.96 8.24 0.90 7.06 0.90
                 7.06 1.12 6.74 1.12 6.74 0.90 4.88 0.90 4.88 1.14 4.56 1.14
                 4.56 0.90 1.20 0.90 1.20 1.62 0.88 1.62 0.88 0.90 0.00 0.90
                 0.00 -0.90 9.60 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  9.60 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 4.66 4.86 4.66 4.62 4.98 4.62 4.98 4.86 6.74 4.86
                 6.74 4.62 7.06 4.62 7.06 4.86 9.60 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  8.12 4.54 7.80 4.54 7.80 4.10 7.54 4.10 7.54 3.74 7.44 3.74
                 7.44 3.42 7.54 3.42 7.54 1.54 7.44 1.54 7.44 1.22 7.86 1.22
                 7.86 3.78 8.12 3.78 ;
        POLYGON  7.22 3.18 7.00 3.18 7.00 4.30 4.66 4.30 4.66 3.90 2.80 3.90
                 2.80 4.54 2.48 4.54 2.48 1.30 2.80 1.30 2.80 3.58 4.98 3.58
                 4.98 3.98 6.68 3.98 6.68 2.86 7.22 2.86 ;
        POLYGON  6.36 1.54 6.32 1.54 6.32 1.80 5.97 2.15 5.97 2.71 6.32 3.06
                 6.32 3.34 6.36 3.34 6.36 3.66 6.00 3.66 6.00 3.20 5.65 2.85
                 5.65 2.01 6.00 1.66 6.00 1.22 6.36 1.22 ;
        POLYGON  5.68 3.66 5.36 3.66 5.36 3.48 5.14 3.26 4.66 3.26 4.66 2.58
                 3.70 2.58 3.70 2.26 4.66 2.26 4.66 1.90 5.26 1.30 5.58 1.30
                 5.58 1.62 5.40 1.62 4.98 2.04 4.98 2.94 5.28 2.94 5.68 3.34 ;
        RECT  3.18 4.22 4.28 4.54 ;
        RECT  3.18 1.58 4.18 1.90 ;
        POLYGON  2.00 2.26 0.18 2.26 0.18 1.30 0.50 1.30 0.50 1.94 1.68 1.94
                 1.68 1.30 2.00 1.30 ;
        POLYGON  1.88 4.54 1.56 4.54 1.56 3.76 0.50 3.76 0.50 4.54 0.18 4.54
                 0.18 3.44 1.88 3.44 ;
    END
END latpq_2

MACRO latpq_1
    CLASS CORE ;
    FOREIGN latpq_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.60 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.08 7.16 2.54 ;
        END
    END gb
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.44 2.40 9.26 2.40 9.26 4.54 8.94 4.54 8.94 1.22 9.26 1.22
                 9.26 2.08 9.44 2.08 ;
        END
    END q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  9.60 0.90 8.56 0.90 8.56 1.54 8.24 1.54 8.24 0.90 7.06 0.90
                 7.06 1.12 6.74 1.12 6.74 0.90 4.88 0.90 4.88 1.14 4.56 1.14
                 4.56 0.90 1.20 0.90 1.20 1.62 0.88 1.62 0.88 0.90 0.00 0.90
                 0.00 -0.90 9.60 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  9.60 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 4.66 4.86 4.66 4.62 4.98 4.62 4.98 4.86 6.74 4.86
                 6.74 4.62 7.06 4.62 7.06 4.86 9.60 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  8.12 4.54 7.80 4.54 7.80 4.10 7.54 4.10 7.54 3.74 7.44 3.74
                 7.44 3.42 7.54 3.42 7.54 1.54 7.44 1.54 7.44 1.22 7.86 1.22
                 7.86 3.78 8.12 3.78 ;
        POLYGON  7.22 3.18 7.00 3.18 7.00 4.30 4.66 4.30 4.66 3.90 2.80 3.90
                 2.80 4.54 2.48 4.54 2.48 1.30 2.80 1.30 2.80 3.58 4.98 3.58
                 4.98 3.98 6.68 3.98 6.68 2.86 7.22 2.86 ;
        POLYGON  6.36 1.54 6.32 1.54 6.32 1.80 5.97 2.15 5.97 2.71 6.32 3.06
                 6.32 3.34 6.36 3.34 6.36 3.66 6.00 3.66 6.00 3.20 5.65 2.85
                 5.65 2.01 6.00 1.66 6.00 1.22 6.36 1.22 ;
        POLYGON  5.68 3.66 5.36 3.66 5.36 3.48 5.14 3.26 4.66 3.26 4.66 2.58
                 3.70 2.58 3.70 2.26 4.66 2.26 4.66 1.90 5.26 1.30 5.58 1.30
                 5.58 1.62 5.40 1.62 4.98 2.04 4.98 2.94 5.28 2.94 5.68 3.34 ;
        RECT  3.18 4.22 4.28 4.54 ;
        RECT  3.18 1.58 4.18 1.90 ;
        POLYGON  2.00 2.26 0.18 2.26 0.18 1.30 0.50 1.30 0.50 1.94 1.68 1.94
                 1.68 1.30 2.00 1.30 ;
        POLYGON  1.88 4.54 1.56 4.54 1.56 3.76 0.50 3.76 0.50 4.54 0.18 4.54
                 0.18 3.44 1.88 3.44 ;
    END
END latpq_1

MACRO latp_4
    CLASS CORE ;
    FOREIGN latp_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.80 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.08 7.12 2.54 ;
        END
    END gb
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.37 3.25 8.60 3.25 8.60 2.93 9.76 2.93 9.76 2.72 10.05 2.72
                 10.05 1.62 8.12 1.62 8.12 1.30 10.37 1.30 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.64 4.53 10.69 4.53 10.69 4.21 12.32 4.21 12.32 1.90
                 10.69 1.90 10.69 1.58 12.64 1.58 ;
        END
    END qb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  12.80 0.90 11.71 0.90 11.71 1.23 11.39 1.23 11.39 0.90
                 7.06 0.90 7.06 1.12 6.74 1.12 6.74 0.90 4.88 0.90 4.88 1.14
                 4.56 1.14 4.56 0.90 1.20 0.90 1.20 1.62 0.88 1.62 0.88 0.90
                 0.00 0.90 0.00 -0.90 12.80 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  12.80 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 4.66 4.86 4.66 4.62 4.98 4.62 4.98 4.86 6.74 4.86
                 6.74 4.62 7.06 4.62 7.06 4.86 9.24 4.86 9.24 4.79 9.66 4.79
                 9.66 4.86 12.80 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  11.71 3.89 9.36 3.89 9.36 4.10 8.12 4.10 8.12 4.54 7.80 4.54
                 7.80 4.10 7.54 4.10 7.54 3.74 7.44 3.74 7.44 3.42 7.54 3.42
                 7.54 2.11 7.44 2.11 7.44 1.22 7.76 1.22 7.76 1.83 7.86 1.83
                 7.86 3.78 9.04 3.78 9.04 3.57 11.39 3.57 11.39 2.34 11.71 2.34 ;
        POLYGON  7.22 3.18 7.00 3.18 7.00 4.30 4.66 4.30 4.66 3.90 2.80 3.90
                 2.80 4.54 2.48 4.54 2.48 1.30 2.80 1.30 2.80 3.58 4.98 3.58
                 4.98 3.98 6.68 3.98 6.68 2.86 7.22 2.86 ;
        POLYGON  6.36 1.54 6.32 1.54 6.32 1.80 5.97 2.15 5.97 2.71 6.32 3.06
                 6.32 3.34 6.36 3.34 6.36 3.66 6.00 3.66 6.00 3.20 5.65 2.85
                 5.65 2.01 6.00 1.66 6.00 1.22 6.36 1.22 ;
        POLYGON  5.68 3.66 5.36 3.66 5.36 3.48 5.14 3.26 4.66 3.26 4.66 2.58
                 3.70 2.58 3.70 2.26 4.66 2.26 4.66 1.90 5.26 1.30 5.58 1.30
                 5.58 1.62 5.40 1.62 4.98 2.04 4.98 2.94 5.28 2.94 5.68 3.34 ;
        RECT  3.18 4.22 4.28 4.54 ;
        RECT  3.18 1.58 4.18 1.90 ;
        POLYGON  2.00 2.26 0.18 2.26 0.18 1.30 0.50 1.30 0.50 1.94 1.68 1.94
                 1.68 1.30 2.00 1.30 ;
        POLYGON  1.88 4.54 1.56 4.54 1.56 3.76 0.50 3.76 0.50 4.54 0.18 4.54
                 0.18 3.44 1.88 3.44 ;
    END
END latp_4

MACRO latp_2
    CLASS CORE ;
    FOREIGN latp_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.24 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.08 7.16 2.54 ;
        END
    END gb
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.73  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.80 1.76 8.50 1.76 8.50 3.46 8.18 3.46 8.18 1.40 8.80 1.40 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.08 4.54 9.66 4.54 9.66 4.22 9.76 4.22 9.76 1.96 9.66 1.96
                 9.66 1.64 10.08 1.64 ;
        END
    END qb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  10.24 0.90 9.28 0.90 9.28 1.08 8.96 1.08 8.96 0.90 7.06 0.90
                 7.06 1.12 6.74 1.12 6.74 0.90 4.88 0.90 4.88 1.14 4.56 1.14
                 4.56 0.90 1.20 0.90 1.20 1.62 0.88 1.62 0.88 0.90 0.00 0.90
                 0.00 -0.90 10.24 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  10.24 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 4.66 4.86 4.66 4.62 4.98 4.62 4.98 4.86 6.74 4.86
                 6.74 4.62 7.06 4.62 7.06 4.86 10.24 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  9.44 2.62 9.34 2.62 9.34 4.10 8.12 4.10 8.12 4.54 7.80 4.54
                 7.80 4.10 7.54 4.10 7.54 3.74 7.44 3.74 7.44 3.42 7.54 3.42
                 7.54 1.54 7.44 1.54 7.44 1.22 7.86 1.22 7.86 3.78 9.02 3.78
                 9.02 2.30 9.44 2.30 ;
        POLYGON  7.22 3.18 7.00 3.18 7.00 4.30 4.66 4.30 4.66 3.90 2.80 3.90
                 2.80 4.54 2.48 4.54 2.48 1.30 2.80 1.30 2.80 3.58 4.98 3.58
                 4.98 3.98 6.68 3.98 6.68 2.86 7.22 2.86 ;
        POLYGON  6.36 1.54 6.32 1.54 6.32 1.80 5.97 2.15 5.97 2.71 6.32 3.06
                 6.32 3.34 6.36 3.34 6.36 3.66 6.00 3.66 6.00 3.20 5.65 2.85
                 5.65 2.01 6.00 1.66 6.00 1.22 6.36 1.22 ;
        POLYGON  5.68 3.66 5.36 3.66 5.36 3.48 5.14 3.26 4.66 3.26 4.66 2.58
                 3.70 2.58 3.70 2.26 4.66 2.26 4.66 1.90 5.26 1.30 5.58 1.30
                 5.58 1.62 5.40 1.62 4.98 2.04 4.98 2.94 5.28 2.94 5.68 3.34 ;
        RECT  3.18 4.22 4.28 4.54 ;
        RECT  3.18 1.58 4.18 1.90 ;
        POLYGON  2.00 2.26 0.18 2.26 0.18 1.30 0.50 1.30 0.50 1.94 1.68 1.94
                 1.68 1.30 2.00 1.30 ;
        POLYGON  1.88 4.54 1.56 4.54 1.56 3.76 0.50 3.76 0.50 4.54 0.18 4.54
                 0.18 3.44 1.88 3.44 ;
    END
END latp_2

MACRO latp_1
    CLASS CORE ;
    FOREIGN latp_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.24 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN gb
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.08 7.16 2.54 ;
        END
    END gb
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.42  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.80 1.76 8.50 1.76 8.50 3.46 8.18 3.46 8.18 1.22 8.58 1.22
                 8.58 1.44 8.80 1.44 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.08 4.30 9.66 4.30 9.66 3.98 9.76 3.98 9.76 1.54 9.66 1.54
                 9.66 1.22 10.08 1.22 ;
        END
    END qb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  10.24 0.90 9.28 0.90 9.28 1.08 8.96 1.08 8.96 0.90 7.06 0.90
                 7.06 1.12 6.74 1.12 6.74 0.90 4.88 0.90 4.88 1.14 4.56 1.14
                 4.56 0.90 1.20 0.90 1.20 1.62 0.88 1.62 0.88 0.90 0.00 0.90
                 0.00 -0.90 10.24 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  10.24 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 4.66 4.86 4.66 4.62 4.98 4.62 4.98 4.86 6.74 4.86
                 6.74 4.62 7.06 4.62 7.06 4.86 10.24 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  9.44 2.62 9.34 2.62 9.34 4.10 8.12 4.10 8.12 4.54 7.80 4.54
                 7.80 4.10 7.54 4.10 7.54 3.74 7.44 3.74 7.44 3.42 7.54 3.42
                 7.54 1.54 7.44 1.54 7.44 1.22 7.86 1.22 7.86 3.78 9.02 3.78
                 9.02 2.30 9.44 2.30 ;
        POLYGON  7.22 3.18 7.00 3.18 7.00 4.30 4.66 4.30 4.66 3.90 2.80 3.90
                 2.80 4.54 2.48 4.54 2.48 1.30 2.80 1.30 2.80 3.58 4.98 3.58
                 4.98 3.98 6.68 3.98 6.68 2.86 7.22 2.86 ;
        POLYGON  6.36 1.54 6.32 1.54 6.32 1.80 5.97 2.15 5.97 2.71 6.32 3.06
                 6.32 3.34 6.36 3.34 6.36 3.66 6.00 3.66 6.00 3.20 5.65 2.85
                 5.65 2.01 6.00 1.66 6.00 1.22 6.36 1.22 ;
        POLYGON  5.68 3.66 5.36 3.66 5.36 3.48 5.14 3.26 4.66 3.26 4.66 2.58
                 3.70 2.58 3.70 2.26 4.66 2.26 4.66 1.90 5.26 1.30 5.58 1.30
                 5.58 1.62 5.40 1.62 4.98 2.04 4.98 2.94 5.28 2.94 5.68 3.34 ;
        RECT  3.18 4.22 4.28 4.54 ;
        RECT  3.18 1.58 4.18 1.90 ;
        POLYGON  2.00 2.26 0.18 2.26 0.18 1.30 0.50 1.30 0.50 1.94 1.68 1.94
                 1.68 1.30 2.00 1.30 ;
        POLYGON  1.88 4.54 1.56 4.54 1.56 3.76 0.50 3.76 0.50 4.54 0.18 4.54
                 0.18 3.44 1.88 3.44 ;
    END
END latp_1

MACRO latnsqb_4
    CLASS CORE ;
    FOREIGN latnsqb_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.64 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.00 2.02 11.32 2.02 11.32 1.70 11.68 1.70 11.68 1.44
                 12.00 1.44 ;
        END
    END g
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.48 4.53 14.58 4.53 14.58 4.21 16.16 4.21 16.16 1.90
                 14.58 1.90 14.58 1.58 16.48 1.58 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 1.92 3.04 2.56 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 0.90 15.60 0.90 15.60 1.23 15.28 1.23 15.28 0.90
                 13.42 0.90 13.42 1.51 13.10 1.51 13.10 0.90 11.74 0.90
                 11.74 1.12 11.42 1.12 11.42 0.90 9.56 0.90 9.56 1.51 9.24 1.51
                 9.24 0.90 0.00 0.90 0.00 -0.90 16.64 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.82 2.58 4.82
                 2.58 4.86 2.94 4.86 2.94 4.62 3.26 4.62 3.26 4.86 9.34 4.86
                 9.34 4.16 9.66 4.16 9.66 4.86 11.42 4.86 11.42 4.16 11.74 4.16
                 11.74 4.86 16.64 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  15.60 3.89 14.21 3.89 14.21 4.10 13.08 4.10 13.08 4.54
                 12.76 4.54 12.76 4.10 12.32 4.10 12.32 1.22 12.64 1.22
                 12.64 3.78 13.89 3.78 13.89 3.57 15.28 3.57 15.28 2.34
                 15.60 2.34 ;
        POLYGON  14.12 1.90 14.10 1.90 14.10 3.00 13.78 3.00 13.78 1.58
                 14.12 1.58 ;
        POLYGON  11.90 2.68 11.68 2.68 11.68 3.84 8.79 3.84 8.79 3.90 6.77 3.90
                 6.77 3.84 5.42 3.84 5.42 4.30 5.10 4.30 5.10 3.66 4.82 3.66
                 4.66 3.50 4.65 3.50 4.65 3.49 4.31 3.15 4.31 2.05 4.92 1.44
                 4.92 1.22 5.24 1.22 5.24 1.58 4.63 2.19 4.63 3.01 4.96 3.34
                 5.42 3.34 5.42 3.52 7.09 3.52 7.09 3.58 8.47 3.58 8.47 3.52
                 11.36 3.52 11.36 2.36 11.90 2.36 ;
        POLYGON  11.04 1.54 11.00 1.54 11.00 2.88 11.04 2.88 11.04 3.20
                 10.68 3.20 10.68 2.48 10.56 2.48 10.56 2.16 10.68 2.16
                 10.68 1.22 11.04 1.22 ;
        POLYGON  10.36 3.20 9.92 3.20 9.92 2.62 5.59 2.62 5.59 2.66 4.95 2.66
                 4.95 2.34 5.27 2.34 5.27 2.30 9.92 2.30 9.92 1.30 10.26 1.30
                 10.26 1.62 10.24 1.62 10.24 2.88 10.36 2.88 ;
        POLYGON  8.98 4.54 5.80 4.54 5.80 4.16 6.12 4.16 6.12 4.22 8.98 4.22 ;
        RECT  5.80 1.22 8.86 1.54 ;
        RECT  7.28 2.94 8.28 3.26 ;
        POLYGON  4.72 4.30 2.50 4.30 2.50 4.50 0.50 4.50 0.50 4.54 0.18 4.54
                 0.18 4.18 2.18 4.18 2.18 3.98 4.72 3.98 ;
        RECT  0.18 1.22 4.36 1.54 ;
        POLYGON  4.04 3.66 3.36 3.66 3.36 3.20 1.96 3.20 1.96 2.88 3.36 2.88
                 3.36 1.86 3.68 1.86 3.68 3.34 4.04 3.34 ;
        RECT  0.88 3.54 1.88 3.86 ;
    END
END latnsqb_4

MACRO latnsqb_2
    CLASS CORE ;
    FOREIGN latnsqb_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.00 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.00 2.02 11.32 2.02 11.32 1.70 11.68 1.70 11.68 1.44
                 12.00 1.44 ;
        END
    END g
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  15.84 2.40 15.72 2.40 15.72 4.54 15.28 4.54 15.28 4.22
                 15.40 4.22 15.40 1.54 15.28 1.54 15.28 1.22 15.72 1.22
                 15.72 2.08 15.84 2.08 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 1.92 3.04 2.56 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 0.90 13.42 0.90 13.42 1.14 13.10 1.14 13.10 0.90
                 11.74 0.90 11.74 1.12 11.42 1.12 11.42 0.90 9.56 0.90
                 9.56 1.54 9.24 1.54 9.24 0.90 0.00 0.90 0.00 -0.90 16.00 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.82 2.58 4.82
                 2.58 4.86 2.94 4.86 2.94 4.62 3.26 4.62 3.26 4.86 9.34 4.86
                 9.34 4.16 9.66 4.16 9.66 4.86 11.42 4.86 11.42 4.16 11.74 4.16
                 11.74 4.86 16.00 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  15.06 2.62 14.98 2.62 14.98 4.10 13.08 4.10 13.08 4.54
                 12.76 4.54 12.76 4.10 12.32 4.10 12.32 1.22 12.64 1.22
                 12.64 3.78 14.66 3.78 14.66 2.30 15.06 2.30 ;
        POLYGON  14.12 1.90 14.10 1.90 14.10 3.08 13.78 3.08 13.78 1.58
                 14.12 1.58 ;
        POLYGON  11.90 2.68 11.68 2.68 11.68 3.84 8.79 3.84 8.79 3.90 6.77 3.90
                 6.77 3.84 5.42 3.84 5.42 4.30 5.10 4.30 5.10 3.66 4.82 3.66
                 4.66 3.50 4.65 3.50 4.65 3.49 4.31 3.15 4.31 2.05 4.92 1.44
                 4.92 1.22 5.24 1.22 5.24 1.58 4.63 2.19 4.63 3.01 4.96 3.34
                 5.42 3.34 5.42 3.52 7.09 3.52 7.09 3.58 8.47 3.58 8.47 3.52
                 11.36 3.52 11.36 2.36 11.90 2.36 ;
        POLYGON  11.04 1.54 11.00 1.54 11.00 2.88 11.04 2.88 11.04 3.20
                 10.68 3.20 10.68 2.48 10.56 2.48 10.56 2.16 10.68 2.16
                 10.68 1.22 11.04 1.22 ;
        POLYGON  10.36 3.20 9.92 3.20 9.92 2.62 5.59 2.62 5.59 2.66 4.95 2.66
                 4.95 2.34 5.27 2.34 5.27 2.30 9.92 2.30 9.92 1.26 10.26 1.26
                 10.26 1.58 10.24 1.58 10.24 2.88 10.36 2.88 ;
        POLYGON  8.98 4.54 5.80 4.54 5.80 4.16 6.12 4.16 6.12 4.22 8.98 4.22 ;
        RECT  5.80 1.22 8.86 1.54 ;
        RECT  7.28 2.94 8.28 3.26 ;
        POLYGON  4.72 4.30 2.50 4.30 2.50 4.50 0.50 4.50 0.50 4.54 0.18 4.54
                 0.18 4.18 2.18 4.18 2.18 3.98 4.72 3.98 ;
        RECT  0.18 1.22 4.36 1.54 ;
        POLYGON  4.04 3.66 3.36 3.66 3.36 3.20 1.96 3.20 1.96 2.88 3.36 2.88
                 3.36 1.86 3.68 1.86 3.68 3.34 4.04 3.34 ;
        RECT  0.88 3.54 1.88 3.86 ;
    END
END latnsqb_2

MACRO latnsqb_1
    CLASS CORE ;
    FOREIGN latnsqb_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.00 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.00 2.02 11.32 2.02 11.32 1.70 11.68 1.70 11.68 1.44
                 12.00 1.44 ;
        END
    END g
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  15.84 2.40 15.72 2.40 15.72 4.54 15.28 4.54 15.28 4.22
                 15.40 4.22 15.40 1.54 15.28 1.54 15.28 1.22 15.72 1.22
                 15.72 2.08 15.84 2.08 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 1.92 3.04 2.56 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 0.90 13.42 0.90 13.42 1.14 13.10 1.14 13.10 0.90
                 11.74 0.90 11.74 1.12 11.42 1.12 11.42 0.90 9.56 0.90
                 9.56 1.54 9.24 1.54 9.24 0.90 0.00 0.90 0.00 -0.90 16.00 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.82 2.58 4.82
                 2.58 4.86 2.94 4.86 2.94 4.62 3.26 4.62 3.26 4.86 9.34 4.86
                 9.34 4.16 9.66 4.16 9.66 4.86 11.42 4.86 11.42 4.16 11.74 4.16
                 11.74 4.86 16.00 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  15.06 2.62 14.98 2.62 14.98 4.10 13.08 4.10 13.08 4.54
                 12.76 4.54 12.76 4.10 12.32 4.10 12.32 1.22 12.64 1.22
                 12.64 3.78 14.66 3.78 14.66 2.30 15.06 2.30 ;
        POLYGON  14.12 1.90 14.10 1.90 14.10 3.00 13.78 3.00 13.78 1.58
                 14.12 1.58 ;
        POLYGON  11.90 2.68 11.68 2.68 11.68 3.84 8.79 3.84 8.79 3.90 6.77 3.90
                 6.77 3.84 5.42 3.84 5.42 4.30 5.10 4.30 5.10 3.66 4.82 3.66
                 4.66 3.50 4.65 3.50 4.65 3.49 4.31 3.15 4.31 2.05 4.92 1.44
                 4.92 1.22 5.24 1.22 5.24 1.58 4.63 2.19 4.63 3.01 4.96 3.34
                 5.42 3.34 5.42 3.52 7.09 3.52 7.09 3.58 8.47 3.58 8.47 3.52
                 11.36 3.52 11.36 2.36 11.90 2.36 ;
        POLYGON  11.04 1.54 11.00 1.54 11.00 2.88 11.04 2.88 11.04 3.20
                 10.68 3.20 10.68 2.48 10.56 2.48 10.56 2.16 10.68 2.16
                 10.68 1.22 11.04 1.22 ;
        POLYGON  10.36 3.20 9.92 3.20 9.92 2.62 5.59 2.62 5.59 2.66 4.95 2.66
                 4.95 2.34 5.27 2.34 5.27 2.30 9.92 2.30 9.92 1.26 10.26 1.26
                 10.26 1.58 10.24 1.58 10.24 2.88 10.36 2.88 ;
        POLYGON  8.98 4.54 5.80 4.54 5.80 4.16 6.12 4.16 6.12 4.22 8.98 4.22 ;
        RECT  5.80 1.22 8.86 1.54 ;
        RECT  7.28 2.94 8.28 3.26 ;
        POLYGON  4.72 4.30 2.50 4.30 2.50 4.50 0.50 4.50 0.50 4.54 0.18 4.54
                 0.18 4.18 2.18 4.18 2.18 3.98 4.72 3.98 ;
        RECT  0.18 1.22 4.36 1.54 ;
        POLYGON  4.04 3.66 3.36 3.66 3.36 3.20 1.96 3.20 1.96 2.88 3.36 2.88
                 3.36 1.86 3.68 1.86 3.68 3.34 4.04 3.34 ;
        RECT  0.88 3.54 1.88 3.86 ;
    END
END latnsqb_1

MACRO latnsq_4
    CLASS CORE ;
    FOREIGN latnsq_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.64 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.00 2.02 11.32 2.02 11.32 1.70 11.68 1.70 11.68 1.44
                 12.00 1.44 ;
        END
    END g
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.20 3.04 15.50 3.04 15.50 3.43 15.18 3.43 15.18 2.72
                 15.88 2.72 15.88 1.68 14.48 1.68 14.48 1.36 16.20 1.36 ;
        END
    END q
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 1.92 3.04 2.56 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 0.90 13.42 0.90 13.42 1.51 13.10 1.51 13.10 0.90
                 11.74 0.90 11.74 1.12 11.42 1.12 11.42 0.90 9.56 0.90
                 9.56 1.51 9.24 1.51 9.24 0.90 0.00 0.90 0.00 -0.90 16.64 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.82 2.58 4.82
                 2.58 4.86 2.94 4.86 2.94 4.62 3.26 4.62 3.26 4.86 9.34 4.86
                 9.34 4.16 9.66 4.16 9.66 4.86 11.42 4.86 11.42 4.16 11.74 4.16
                 11.74 4.86 16.64 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  14.12 1.90 14.10 1.90 14.10 3.01 13.78 3.01 13.78 1.58
                 14.12 1.58 ;
        POLYGON  13.08 4.54 12.76 4.54 12.76 4.10 12.32 4.10 12.32 1.22
                 12.64 1.22 12.64 3.78 13.08 3.78 ;
        POLYGON  11.90 2.68 11.68 2.68 11.68 3.84 8.79 3.84 8.79 3.90 6.77 3.90
                 6.77 3.84 5.42 3.84 5.42 4.30 5.10 4.30 5.10 3.66 4.82 3.66
                 4.66 3.50 4.65 3.50 4.65 3.49 4.31 3.15 4.31 2.05 4.92 1.44
                 4.92 1.22 5.24 1.22 5.24 1.58 4.63 2.19 4.63 3.01 4.96 3.34
                 5.42 3.34 5.42 3.52 7.09 3.52 7.09 3.58 8.47 3.58 8.47 3.52
                 11.36 3.52 11.36 2.36 11.90 2.36 ;
        POLYGON  11.04 1.54 11.00 1.54 11.00 2.88 11.04 2.88 11.04 3.20
                 10.68 3.20 10.68 2.48 10.56 2.48 10.56 2.16 10.68 2.16
                 10.68 1.22 11.04 1.22 ;
        POLYGON  10.36 3.20 9.92 3.20 9.92 2.62 5.59 2.62 5.59 2.66 4.95 2.66
                 4.95 2.34 5.27 2.34 5.27 2.30 9.92 2.30 9.92 1.30 10.26 1.30
                 10.26 1.62 10.24 1.62 10.24 2.88 10.36 2.88 ;
        POLYGON  8.98 4.54 5.80 4.54 5.80 4.16 6.12 4.16 6.12 4.22 8.98 4.22 ;
        RECT  5.80 1.22 8.86 1.54 ;
        RECT  7.28 2.94 8.28 3.26 ;
        POLYGON  4.72 4.30 2.50 4.30 2.50 4.50 0.50 4.50 0.50 4.54 0.18 4.54
                 0.18 4.18 2.18 4.18 2.18 3.98 4.72 3.98 ;
        RECT  0.18 1.22 4.36 1.54 ;
        POLYGON  4.04 3.66 3.36 3.66 3.36 3.20 1.96 3.20 1.96 2.88 3.36 2.88
                 3.36 1.86 3.68 1.86 3.68 3.34 4.04 3.34 ;
        RECT  0.88 3.54 1.88 3.86 ;
    END
END latnsq_4

MACRO latnsq_2
    CLASS CORE ;
    FOREIGN latnsq_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.00 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.00 2.02 11.32 2.02 11.32 1.70 11.68 1.70 11.68 1.44
                 12.00 1.44 ;
        END
    END g
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.80  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  15.20 2.40 14.76 2.40 14.76 4.54 14.42 4.54 14.42 3.14
                 14.44 3.14 14.44 1.33 14.80 1.33 14.80 2.08 15.20 2.08 ;
        END
    END q
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 1.92 3.04 2.56 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 0.90 15.50 0.90 15.50 1.20 15.18 1.20 15.18 0.90
                 13.42 0.90 13.42 1.51 13.10 1.51 13.10 0.90 11.74 0.90
                 11.74 1.12 11.42 1.12 11.42 0.90 9.56 0.90 9.56 1.54 9.24 1.54
                 9.24 0.90 0.00 0.90 0.00 -0.90 16.00 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.82 2.58 4.82
                 2.58 4.86 2.94 4.86 2.94 4.62 3.26 4.62 3.26 4.86 9.34 4.86
                 9.34 4.16 9.66 4.16 9.66 4.86 11.42 4.86 11.42 4.16 11.74 4.16
                 11.74 4.86 15.18 4.86 15.18 4.22 15.50 4.22 15.50 4.86
                 16.00 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  14.12 1.90 14.10 1.90 14.10 3.08 13.78 3.08 13.78 1.58
                 14.12 1.58 ;
        POLYGON  13.08 4.54 12.76 4.54 12.76 4.10 12.32 4.10 12.32 1.22
                 12.64 1.22 12.64 3.78 13.08 3.78 ;
        POLYGON  11.90 2.68 11.68 2.68 11.68 3.84 8.79 3.84 8.79 3.90 6.77 3.90
                 6.77 3.84 5.42 3.84 5.42 4.30 5.10 4.30 5.10 3.66 4.82 3.66
                 4.66 3.50 4.65 3.50 4.65 3.49 4.31 3.15 4.31 2.05 4.92 1.44
                 4.92 1.22 5.24 1.22 5.24 1.58 4.63 2.19 4.63 3.01 4.96 3.34
                 5.42 3.34 5.42 3.52 7.09 3.52 7.09 3.58 8.47 3.58 8.47 3.52
                 11.36 3.52 11.36 2.36 11.90 2.36 ;
        POLYGON  11.04 1.54 11.00 1.54 11.00 2.88 11.04 2.88 11.04 3.20
                 10.68 3.20 10.68 2.48 10.56 2.48 10.56 2.16 10.68 2.16
                 10.68 1.22 11.04 1.22 ;
        POLYGON  10.36 3.20 9.92 3.20 9.92 2.62 5.59 2.62 5.59 2.66 4.95 2.66
                 4.95 2.34 5.27 2.34 5.27 2.30 9.92 2.30 9.92 1.22 10.26 1.22
                 10.26 1.54 10.24 1.54 10.24 2.88 10.36 2.88 ;
        POLYGON  8.98 4.54 5.80 4.54 5.80 4.16 6.12 4.16 6.12 4.22 8.98 4.22 ;
        RECT  5.80 1.22 8.86 1.54 ;
        RECT  7.28 2.94 8.28 3.26 ;
        POLYGON  4.72 4.30 2.50 4.30 2.50 4.50 0.50 4.50 0.50 4.54 0.18 4.54
                 0.18 4.18 2.18 4.18 2.18 3.98 4.72 3.98 ;
        RECT  0.18 1.22 4.36 1.54 ;
        POLYGON  4.04 3.66 3.36 3.66 3.36 3.20 1.96 3.20 1.96 2.88 3.36 2.88
                 3.36 1.86 3.68 1.86 3.68 3.34 4.04 3.34 ;
        RECT  0.88 3.54 1.88 3.86 ;
    END
END latnsq_2

MACRO latnsq_1
    CLASS CORE ;
    FOREIGN latnsq_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.00 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.00 2.02 11.32 2.02 11.32 1.70 11.68 1.70 11.68 1.44
                 12.00 1.44 ;
        END
    END g
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.29  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  15.20 2.40 14.76 2.40 14.76 4.25 14.42 4.25 14.42 3.14
                 14.44 3.14 14.44 1.22 14.80 1.22 14.80 2.08 15.20 2.08 ;
        END
    END q
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 1.92 3.04 2.56 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 0.90 15.50 0.90 15.50 1.20 15.18 1.20 15.18 0.90
                 13.42 0.90 13.42 1.51 13.10 1.51 13.10 0.90 11.74 0.90
                 11.74 1.12 11.42 1.12 11.42 0.90 9.56 0.90 9.56 1.50 9.24 1.50
                 9.24 0.90 0.00 0.90 0.00 -0.90 16.00 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.82 2.58 4.82
                 2.58 4.86 2.94 4.86 2.94 4.62 3.26 4.62 3.26 4.86 9.34 4.86
                 9.34 4.16 9.66 4.16 9.66 4.86 11.42 4.86 11.42 4.16 11.74 4.16
                 11.74 4.86 15.18 4.86 15.18 4.22 15.50 4.22 15.50 4.86
                 16.00 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  14.12 1.90 14.10 1.90 14.10 3.08 13.78 3.08 13.78 1.58
                 14.12 1.58 ;
        POLYGON  13.08 4.54 12.76 4.54 12.76 4.10 12.32 4.10 12.32 1.22
                 12.64 1.22 12.64 3.78 13.08 3.78 ;
        POLYGON  11.90 2.68 11.68 2.68 11.68 3.84 8.79 3.84 8.79 3.90 6.77 3.90
                 6.77 3.84 5.42 3.84 5.42 4.30 5.10 4.30 5.10 3.66 4.82 3.66
                 4.66 3.50 4.65 3.50 4.65 3.49 4.31 3.15 4.31 2.05 4.92 1.44
                 4.92 1.22 5.24 1.22 5.24 1.58 4.63 2.19 4.63 3.01 4.96 3.34
                 5.42 3.34 5.42 3.52 7.09 3.52 7.09 3.58 8.47 3.58 8.47 3.52
                 11.36 3.52 11.36 2.36 11.90 2.36 ;
        POLYGON  11.04 1.54 11.00 1.54 11.00 2.88 11.04 2.88 11.04 3.20
                 10.68 3.20 10.68 2.48 10.56 2.48 10.56 2.16 10.68 2.16
                 10.68 1.22 11.04 1.22 ;
        POLYGON  10.36 3.20 9.92 3.20 9.92 2.62 5.59 2.62 5.59 2.66 4.95 2.66
                 4.95 2.34 5.27 2.34 5.27 2.30 9.92 2.30 9.92 1.30 10.26 1.30
                 10.26 1.62 10.24 1.62 10.24 2.88 10.36 2.88 ;
        POLYGON  8.98 4.54 5.80 4.54 5.80 4.16 6.12 4.16 6.12 4.22 8.98 4.22 ;
        RECT  5.80 1.22 8.86 1.54 ;
        RECT  7.28 2.94 8.28 3.26 ;
        POLYGON  4.72 4.30 2.50 4.30 2.50 4.50 0.50 4.50 0.50 4.54 0.18 4.54
                 0.18 4.18 2.18 4.18 2.18 3.98 4.72 3.98 ;
        RECT  0.18 1.22 4.36 1.54 ;
        POLYGON  4.04 3.66 3.36 3.66 3.36 3.20 1.96 3.20 1.96 2.88 3.36 2.88
                 3.36 1.86 3.68 1.86 3.68 3.34 4.04 3.34 ;
        RECT  0.88 3.54 1.88 3.86 ;
    END
END latnsq_1

MACRO latns_4
    CLASS CORE ;
    FOREIGN latns_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.56 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.00 2.02 11.32 2.02 11.32 1.70 11.68 1.70 11.68 1.44
                 12.00 1.44 ;
        END
    END g
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.20 3.04 15.50 3.04 15.50 3.43 15.18 3.43 15.18 2.72
                 15.88 2.72 15.88 1.68 14.48 1.68 14.48 1.36 16.20 1.36 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  18.40 4.53 16.56 4.53 16.56 4.21 18.08 4.21 18.08 1.90
                 16.56 1.90 16.56 1.58 18.40 1.58 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 1.92 3.04 2.56 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  18.56 0.90 17.58 0.90 17.58 1.23 17.26 1.23 17.26 0.90
                 13.42 0.90 13.42 1.51 13.10 1.51 13.10 0.90 11.74 0.90
                 11.74 1.12 11.42 1.12 11.42 0.90 9.56 0.90 9.56 1.51 9.24 1.51
                 9.24 0.90 0.00 0.90 0.00 -0.90 18.56 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  18.56 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.82 2.58 4.82
                 2.58 4.86 2.94 4.86 2.94 4.62 3.26 4.62 3.26 4.86 9.34 4.86
                 9.34 4.16 9.66 4.16 9.66 4.86 11.42 4.86 11.42 4.16 11.74 4.16
                 11.74 4.86 18.56 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  17.58 3.89 16.19 3.89 16.19 4.10 13.08 4.10 13.08 4.54
                 12.76 4.54 12.76 4.10 12.32 4.10 12.32 1.22 12.64 1.22
                 12.64 3.78 15.87 3.78 15.87 3.57 17.26 3.57 17.26 2.34
                 17.58 2.34 ;
        POLYGON  14.12 1.90 14.10 1.90 14.10 3.01 13.78 3.01 13.78 1.58
                 14.12 1.58 ;
        POLYGON  11.90 2.68 11.68 2.68 11.68 3.84 8.79 3.84 8.79 3.90 6.77 3.90
                 6.77 3.84 5.42 3.84 5.42 4.30 5.10 4.30 5.10 3.66 4.82 3.66
                 4.66 3.50 4.65 3.50 4.65 3.49 4.31 3.15 4.31 2.05 4.92 1.44
                 4.92 1.22 5.24 1.22 5.24 1.58 4.63 2.19 4.63 3.01 4.96 3.34
                 5.42 3.34 5.42 3.52 7.09 3.52 7.09 3.58 8.47 3.58 8.47 3.52
                 11.36 3.52 11.36 2.36 11.90 2.36 ;
        POLYGON  11.04 1.54 11.00 1.54 11.00 2.88 11.04 2.88 11.04 3.20
                 10.68 3.20 10.68 2.48 10.56 2.48 10.56 2.16 10.68 2.16
                 10.68 1.22 11.04 1.22 ;
        POLYGON  10.36 3.20 9.92 3.20 9.92 2.62 5.59 2.62 5.59 2.66 4.95 2.66
                 4.95 2.34 5.27 2.34 5.27 2.30 9.92 2.30 9.92 1.30 10.26 1.30
                 10.26 1.62 10.24 1.62 10.24 2.88 10.36 2.88 ;
        POLYGON  8.98 4.54 5.80 4.54 5.80 4.16 6.12 4.16 6.12 4.22 8.98 4.22 ;
        RECT  5.80 1.22 8.86 1.54 ;
        RECT  7.28 2.94 8.28 3.26 ;
        POLYGON  4.72 4.30 2.50 4.30 2.50 4.50 0.50 4.50 0.50 4.54 0.18 4.54
                 0.18 4.18 2.18 4.18 2.18 3.98 4.72 3.98 ;
        RECT  0.18 1.22 4.36 1.54 ;
        POLYGON  4.04 3.66 3.36 3.66 3.36 3.20 1.96 3.20 1.96 2.88 3.36 2.88
                 3.36 1.86 3.68 1.86 3.68 3.34 4.04 3.34 ;
        RECT  0.88 3.54 1.88 3.86 ;
    END
END latns_4

MACRO latns_2
    CLASS CORE ;
    FOREIGN latns_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.64 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.00 2.02 11.32 2.02 11.32 1.70 11.68 1.70 11.68 1.44
                 12.00 1.44 ;
        END
    END g
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.74  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  15.20 1.76 14.76 1.76 14.76 3.46 14.40 3.46 14.40 3.14
                 14.44 3.14 14.44 1.22 14.80 1.22 14.80 1.44 15.20 1.44 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.48 2.40 16.32 2.40 16.32 4.54 15.88 4.54 15.88 4.22
                 16.00 4.22 16.00 1.54 15.88 1.54 15.88 1.22 16.32 1.22
                 16.32 2.08 16.48 2.08 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 1.92 3.04 2.56 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 0.90 13.42 0.90 13.42 1.52 13.10 1.52 13.10 0.90
                 11.74 0.90 11.74 1.12 11.42 1.12 11.42 0.90 9.56 0.90
                 9.56 1.54 9.24 1.54 9.24 0.90 0.00 0.90 0.00 -0.90 16.64 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.82 2.58 4.82
                 2.58 4.86 2.94 4.86 2.94 4.62 3.26 4.62 3.26 4.86 9.34 4.86
                 9.34 4.16 9.66 4.16 9.66 4.86 11.42 4.86 11.42 4.16 11.74 4.16
                 11.74 4.86 16.64 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  15.66 2.62 15.58 2.62 15.58 4.10 13.08 4.10 13.08 4.54
                 12.76 4.54 12.76 4.10 12.32 4.10 12.32 1.22 12.64 1.22
                 12.64 3.78 15.26 3.78 15.26 2.30 15.66 2.30 ;
        POLYGON  14.12 1.90 14.10 1.90 14.10 3.00 13.78 3.00 13.78 1.58
                 14.12 1.58 ;
        POLYGON  11.90 2.68 11.68 2.68 11.68 3.84 8.79 3.84 8.79 3.90 6.77 3.90
                 6.77 3.84 5.42 3.84 5.42 4.30 5.10 4.30 5.10 3.66 4.82 3.66
                 4.66 3.50 4.65 3.50 4.65 3.49 4.31 3.15 4.31 2.05 4.92 1.44
                 4.92 1.22 5.24 1.22 5.24 1.58 4.63 2.19 4.63 3.01 4.96 3.34
                 5.42 3.34 5.42 3.52 7.09 3.52 7.09 3.58 8.47 3.58 8.47 3.52
                 11.36 3.52 11.36 2.36 11.90 2.36 ;
        POLYGON  11.04 1.54 11.00 1.54 11.00 2.88 11.04 2.88 11.04 3.20
                 10.68 3.20 10.68 2.48 10.56 2.48 10.56 2.16 10.68 2.16
                 10.68 1.22 11.04 1.22 ;
        POLYGON  10.36 3.20 9.92 3.20 9.92 2.62 5.59 2.62 5.59 2.66 4.95 2.66
                 4.95 2.34 5.27 2.34 5.27 2.30 9.92 2.30 9.92 1.26 10.26 1.26
                 10.26 1.58 10.24 1.58 10.24 2.88 10.36 2.88 ;
        POLYGON  8.98 4.54 5.80 4.54 5.80 4.16 6.12 4.16 6.12 4.22 8.98 4.22 ;
        RECT  5.80 1.22 8.86 1.54 ;
        RECT  7.28 2.94 8.28 3.26 ;
        POLYGON  4.72 4.30 2.50 4.30 2.50 4.50 0.50 4.50 0.50 4.54 0.18 4.54
                 0.18 4.18 2.18 4.18 2.18 3.98 4.72 3.98 ;
        RECT  0.18 1.22 4.36 1.54 ;
        POLYGON  4.04 3.66 3.36 3.66 3.36 3.20 1.96 3.20 1.96 2.88 3.36 2.88
                 3.36 1.86 3.68 1.86 3.68 3.34 4.04 3.34 ;
        RECT  0.88 3.54 1.88 3.86 ;
    END
END latns_2

MACRO latns_1
    CLASS CORE ;
    FOREIGN latns_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.64 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.00 2.02 11.32 2.02 11.32 1.70 11.68 1.70 11.68 1.44
                 12.00 1.44 ;
        END
    END g
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.39  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  15.20 1.76 14.76 1.76 14.76 3.46 14.40 3.46 14.40 3.14
                 14.44 3.14 14.44 1.22 14.80 1.22 14.80 1.44 15.20 1.44 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.48 2.40 16.32 2.40 16.32 4.54 15.88 4.54 15.88 4.22
                 16.00 4.22 16.00 1.54 15.88 1.54 15.88 1.22 16.32 1.22
                 16.32 2.08 16.48 2.08 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 1.92 3.04 2.56 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 0.90 13.42 0.90 13.42 1.14 13.10 1.14 13.10 0.90
                 11.74 0.90 11.74 1.12 11.42 1.12 11.42 0.90 9.56 0.90
                 9.56 1.54 9.24 1.54 9.24 0.90 0.00 0.90 0.00 -0.90 16.64 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.82 2.58 4.82
                 2.58 4.86 2.94 4.86 2.94 4.62 3.26 4.62 3.26 4.86 9.34 4.86
                 9.34 4.16 9.66 4.16 9.66 4.86 11.42 4.86 11.42 4.16 11.74 4.16
                 11.74 4.86 16.64 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  15.66 2.62 15.58 2.62 15.58 4.10 13.08 4.10 13.08 4.54
                 12.76 4.54 12.76 4.10 12.32 4.10 12.32 1.22 12.64 1.22
                 12.64 3.78 15.26 3.78 15.26 2.30 15.66 2.30 ;
        POLYGON  14.12 1.90 14.10 1.90 14.10 3.00 13.78 3.00 13.78 1.58
                 14.12 1.58 ;
        POLYGON  11.90 2.68 11.68 2.68 11.68 3.84 8.79 3.84 8.79 3.90 6.77 3.90
                 6.77 3.84 5.42 3.84 5.42 4.30 5.10 4.30 5.10 3.66 4.82 3.66
                 4.66 3.50 4.65 3.50 4.65 3.49 4.31 3.15 4.31 2.05 4.92 1.44
                 4.92 1.22 5.24 1.22 5.24 1.58 4.63 2.19 4.63 3.01 4.96 3.34
                 5.42 3.34 5.42 3.52 7.09 3.52 7.09 3.58 8.47 3.58 8.47 3.52
                 11.36 3.52 11.36 2.36 11.90 2.36 ;
        POLYGON  11.04 1.54 11.00 1.54 11.00 2.88 11.04 2.88 11.04 3.20
                 10.68 3.20 10.68 2.48 10.56 2.48 10.56 2.16 10.68 2.16
                 10.68 1.22 11.04 1.22 ;
        POLYGON  10.36 3.20 9.92 3.20 9.92 2.62 5.59 2.62 5.59 2.66 4.95 2.66
                 4.95 2.34 5.27 2.34 5.27 2.30 9.92 2.30 9.92 1.26 10.26 1.26
                 10.26 1.58 10.24 1.58 10.24 2.88 10.36 2.88 ;
        POLYGON  8.98 4.54 5.80 4.54 5.80 4.16 6.12 4.16 6.12 4.22 8.98 4.22 ;
        RECT  5.80 1.22 8.86 1.54 ;
        RECT  7.28 2.94 8.28 3.26 ;
        POLYGON  4.72 4.30 2.50 4.30 2.50 4.50 0.50 4.50 0.50 4.54 0.18 4.54
                 0.18 4.18 2.18 4.18 2.18 3.98 4.72 3.98 ;
        RECT  0.18 1.22 4.36 1.54 ;
        POLYGON  4.04 3.66 3.36 3.66 3.36 3.20 1.96 3.20 1.96 2.88 3.36 2.88
                 3.36 1.86 3.68 1.86 3.68 3.34 4.04 3.34 ;
        RECT  0.88 3.54 1.88 3.86 ;
    END
END latns_1

MACRO latnrsqb_4
    CLASS CORE ;
    FOREIGN latnrsqb_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.76 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.24 2.72 3.68 3.22 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.58 2.72 14.26 2.72 14.26 2.40 14.24 2.40 14.24 2.08
                 14.58 2.08 ;
        END
    END g
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  21.60 4.53 19.41 4.53 19.41 4.21 21.28 4.21 21.28 1.90
                 19.41 1.90 19.41 1.58 21.60 1.58 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  18.08 1.22 18.59 1.86 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.90  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.71 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.76 0.90 20.43 0.90 20.43 1.23 20.11 1.23 20.11 0.90
                 17.69 0.90 17.69 1.28 17.37 1.28 17.37 0.90 14.78 0.90
                 14.78 1.50 14.46 1.50 14.46 0.90 12.60 0.90 12.60 1.28
                 12.28 1.28 12.28 0.90 8.24 0.90 8.24 1.24 7.92 1.24 7.92 0.90
                 1.20 0.90 1.20 1.28 0.88 1.28 0.88 0.90 0.00 0.90 0.00 -0.90
                 21.76 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.76 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.16 1.20 4.16
                 1.20 4.86 1.56 4.86 1.56 4.16 1.88 4.16 1.88 4.86 12.28 4.86
                 12.28 4.16 12.60 4.16 12.60 4.86 14.42 4.86 14.42 4.16
                 15.30 4.16 15.30 4.86 16.67 4.86 16.67 2.95 16.99 2.95
                 16.99 4.86 21.76 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.43 3.89 19.09 3.89 19.09 4.54 17.43 4.54 17.43 2.52
                 16.21 2.52 16.21 3.84 15.89 3.84 15.89 2.18 15.46 2.18
                 15.28 2.00 15.28 1.22 15.60 1.22 15.60 1.86 16.21 1.86
                 16.21 2.20 17.75 2.20 17.75 4.22 18.77 4.22 18.77 3.57
                 20.11 3.57 20.11 2.34 20.43 2.34 ;
        RECT  18.73 2.23 19.05 3.25 ;
        RECT  15.98 1.22 16.99 1.54 ;
        POLYGON  15.22 3.84 5.34 3.84 5.34 4.30 5.02 4.30 5.02 3.84 4.70 3.84
                 4.70 1.90 5.02 1.90 5.02 3.52 14.90 3.52 14.90 2.40 15.22 2.40 ;
        POLYGON  14.08 1.54 13.94 1.54 13.94 1.95 13.82 2.07 13.82 2.48
                 13.94 2.60 13.94 2.88 13.98 2.88 13.98 3.20 13.62 3.20
                 13.62 2.74 13.50 2.62 13.50 1.93 13.62 1.81 13.62 1.22
                 14.08 1.22 ;
        POLYGON  13.30 1.62 13.18 1.74 13.18 2.88 13.30 2.88 13.30 3.20
                 5.34 3.20 5.34 2.44 5.66 2.44 5.66 2.88 12.86 2.88 12.86 1.47
                 12.91 1.47 12.91 1.37 12.98 1.37 12.98 1.30 13.30 1.30 ;
        POLYGON  11.92 1.60 11.60 1.60 11.60 1.54 8.88 1.54 8.88 1.88 7.28 1.88
                 7.28 1.60 6.46 1.60 6.46 1.28 7.60 1.28 7.60 1.56 8.56 1.56
                 8.56 1.22 11.92 1.22 ;
        POLYGON  11.92 4.54 5.72 4.54 5.72 4.16 6.04 4.16 6.04 4.22 11.92 4.22 ;
        POLYGON  11.22 2.52 8.70 2.52 8.70 2.20 10.90 2.20 10.90 2.04
                 11.22 2.04 ;
        POLYGON  7.46 2.52 6.46 2.52 5.82 1.88 5.82 1.54 4.38 1.54 4.38 2.24
                 2.04 2.24 2.04 1.22 2.36 1.22 2.36 1.92 4.06 1.92 4.06 1.22
                 6.14 1.22 6.14 1.74 6.60 2.20 7.46 2.20 ;
        POLYGON  4.64 4.50 3.96 4.50 3.96 4.54 3.64 4.54 3.64 4.18 4.64 4.18 ;
        POLYGON  3.74 1.60 3.42 1.60 3.42 1.54 2.74 1.54 2.74 1.22 3.74 1.22 ;
        RECT  2.26 4.22 3.26 4.54 ;
        POLYGON  2.18 3.42 0.50 3.42 0.50 4.48 0.16 4.48 0.16 1.22 0.50 1.22
                 0.50 1.54 0.48 1.54 0.48 3.10 2.18 3.10 ;
    END
END latnrsqb_4

MACRO latnrsqb_2
    CLASS CORE ;
    FOREIGN latnrsqb_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.24 2.72 3.68 3.22 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.58 2.72 14.26 2.72 14.26 2.40 14.24 2.40 14.24 2.08
                 14.58 2.08 ;
        END
    END g
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.71  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.96 2.40 20.47 2.40 20.47 4.54 20.13 4.54 20.13 4.22
                 20.15 4.22 20.15 1.80 20.03 1.80 20.03 1.48 20.47 1.48
                 20.47 2.08 20.96 2.08 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  18.08 1.22 18.59 1.86 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.90  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.71 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 0.90 19.65 0.90 19.65 1.92 19.33 1.92 19.33 0.90
                 17.69 0.90 17.69 1.28 17.37 1.28 17.37 0.90 14.78 0.90
                 14.78 1.14 14.46 1.14 14.46 0.90 12.60 0.90 12.60 1.28
                 12.28 1.28 12.28 0.90 8.24 0.90 8.24 1.24 7.92 1.24 7.92 0.90
                 1.20 0.90 1.20 1.58 0.88 1.58 0.88 0.90 0.00 0.90 0.00 -0.90
                 21.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.16 1.20 4.16
                 1.20 4.86 1.56 4.86 1.56 4.16 1.88 4.16 1.88 4.86 12.28 4.86
                 12.28 4.16 12.60 4.16 12.60 4.86 14.42 4.86 14.42 4.16
                 15.30 4.16 15.30 4.86 16.67 4.86 16.67 2.95 16.99 2.95
                 16.99 4.86 21.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  19.81 4.54 17.43 4.54 17.43 2.52 16.21 2.52 16.21 3.84
                 15.89 3.84 15.89 2.18 15.46 2.18 15.28 2.00 15.28 1.22
                 15.60 1.22 15.60 1.86 16.21 1.86 16.21 2.20 17.75 2.20
                 17.75 4.22 19.49 4.22 19.49 2.28 19.81 2.28 ;
        RECT  18.73 2.76 19.05 3.90 ;
        RECT  15.98 1.22 16.99 1.54 ;
        POLYGON  15.22 3.84 5.34 3.84 5.34 4.30 5.02 4.30 5.02 3.84 4.70 3.84
                 4.70 1.90 5.02 1.90 5.02 3.52 14.90 3.52 14.90 2.40 15.22 2.40 ;
        POLYGON  14.08 1.54 13.94 1.54 13.94 1.95 13.82 2.07 13.82 2.48
                 13.94 2.60 13.94 2.88 13.98 2.88 13.98 3.20 13.62 3.20
                 13.62 2.74 13.50 2.62 13.50 1.93 13.62 1.81 13.62 1.22
                 14.08 1.22 ;
        POLYGON  13.30 1.62 13.18 1.74 13.18 2.88 13.30 2.88 13.30 3.20
                 5.34 3.20 5.34 2.44 5.66 2.44 5.66 2.88 12.86 2.88 12.86 1.47
                 12.91 1.47 12.91 1.37 12.98 1.37 12.98 1.30 13.30 1.30 ;
        POLYGON  11.92 1.60 11.60 1.60 11.60 1.54 8.88 1.54 8.88 1.88 7.28 1.88
                 7.28 1.60 6.46 1.60 6.46 1.28 7.60 1.28 7.60 1.56 8.56 1.56
                 8.56 1.22 11.92 1.22 ;
        POLYGON  11.92 4.54 5.72 4.54 5.72 4.16 6.04 4.16 6.04 4.22 11.92 4.22 ;
        POLYGON  11.22 2.52 8.70 2.52 8.70 2.20 10.90 2.20 10.90 2.04
                 11.22 2.04 ;
        POLYGON  7.46 2.52 6.46 2.52 5.82 1.88 5.82 1.54 4.38 1.54 4.38 2.24
                 2.04 2.24 2.04 1.22 2.36 1.22 2.36 1.92 4.06 1.92 4.06 1.22
                 6.14 1.22 6.14 1.74 6.60 2.20 7.46 2.20 ;
        POLYGON  4.64 4.50 3.96 4.50 3.96 4.54 3.64 4.54 3.64 4.18 4.64 4.18 ;
        POLYGON  3.74 1.60 3.42 1.60 3.42 1.54 2.74 1.54 2.74 1.22 3.74 1.22 ;
        RECT  2.26 4.22 3.26 4.54 ;
        POLYGON  2.18 3.42 0.50 3.42 0.50 4.48 0.16 4.48 0.16 1.22 0.50 1.22
                 0.50 1.54 0.48 1.54 0.48 3.10 2.18 3.10 ;
    END
END latnrsqb_2

MACRO latnrsqb_1
    CLASS CORE ;
    FOREIGN latnrsqb_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.24 2.72 3.68 3.22 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.58 2.72 14.26 2.72 14.26 2.40 14.24 2.40 14.24 2.08
                 14.58 2.08 ;
        END
    END g
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.23  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.96 2.40 20.47 2.40 20.47 4.54 20.13 4.54 20.13 4.22
                 20.15 4.22 20.15 1.54 20.03 1.54 20.03 1.22 20.47 1.22
                 20.47 2.08 20.96 2.08 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  18.08 1.22 18.59 1.86 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.90  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.71 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 0.90 19.65 0.90 19.65 1.66 19.33 1.66 19.33 0.90
                 17.69 0.90 17.69 1.28 17.37 1.28 17.37 0.90 14.78 0.90
                 14.78 1.14 14.46 1.14 14.46 0.90 12.60 0.90 12.60 1.28
                 12.28 1.28 12.28 0.90 8.24 0.90 8.24 1.24 7.92 1.24 7.92 0.90
                 1.20 0.90 1.20 1.58 0.88 1.58 0.88 0.90 0.00 0.90 0.00 -0.90
                 21.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.16 1.20 4.16
                 1.20 4.86 1.56 4.86 1.56 4.16 1.88 4.16 1.88 4.86 12.28 4.86
                 12.28 4.16 12.60 4.16 12.60 4.86 14.42 4.86 14.42 4.16
                 15.30 4.16 15.30 4.86 16.67 4.86 16.67 2.95 16.99 2.95
                 16.99 4.86 21.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  19.81 4.54 17.43 4.54 17.43 2.52 16.21 2.52 16.21 3.84
                 15.89 3.84 15.89 2.18 15.46 2.18 15.28 2.00 15.28 1.22
                 15.60 1.22 15.60 1.86 16.21 1.86 16.21 2.20 17.75 2.20
                 17.75 4.22 19.49 4.22 19.49 2.28 19.81 2.28 ;
        RECT  18.73 2.76 19.05 3.90 ;
        RECT  15.98 1.22 16.99 1.54 ;
        POLYGON  15.22 3.84 5.34 3.84 5.34 4.30 5.02 4.30 5.02 3.84 4.70 3.84
                 4.70 1.90 5.02 1.90 5.02 3.52 14.90 3.52 14.90 2.40 15.22 2.40 ;
        POLYGON  14.08 1.54 13.94 1.54 13.94 1.95 13.82 2.07 13.82 2.48
                 13.94 2.60 13.94 2.88 13.98 2.88 13.98 3.20 13.62 3.20
                 13.62 2.74 13.50 2.62 13.50 1.93 13.62 1.81 13.62 1.22
                 14.08 1.22 ;
        POLYGON  13.30 1.62 13.18 1.74 13.18 2.88 13.30 2.88 13.30 3.20
                 5.34 3.20 5.34 2.44 5.66 2.44 5.66 2.88 12.86 2.88 12.86 1.47
                 12.91 1.47 12.91 1.37 12.98 1.37 12.98 1.30 13.30 1.30 ;
        POLYGON  11.92 1.60 11.60 1.60 11.60 1.54 8.88 1.54 8.88 1.88 7.28 1.88
                 7.28 1.60 6.46 1.60 6.46 1.28 7.60 1.28 7.60 1.56 8.56 1.56
                 8.56 1.22 11.92 1.22 ;
        POLYGON  11.92 4.54 5.72 4.54 5.72 4.16 6.04 4.16 6.04 4.22 11.92 4.22 ;
        POLYGON  11.22 2.52 8.70 2.52 8.70 2.20 10.90 2.20 10.90 2.04
                 11.22 2.04 ;
        POLYGON  7.46 2.52 6.46 2.52 5.82 1.88 5.82 1.54 4.38 1.54 4.38 2.24
                 2.04 2.24 2.04 1.22 2.36 1.22 2.36 1.92 4.06 1.92 4.06 1.22
                 6.14 1.22 6.14 1.74 6.60 2.20 7.46 2.20 ;
        POLYGON  4.64 4.50 3.96 4.50 3.96 4.54 3.64 4.54 3.64 4.18 4.64 4.18 ;
        POLYGON  3.74 1.60 3.42 1.60 3.42 1.54 2.74 1.54 2.74 1.22 3.74 1.22 ;
        RECT  2.26 4.22 3.26 4.54 ;
        POLYGON  2.18 3.42 0.50 3.42 0.50 4.48 0.16 4.48 0.16 1.22 0.50 1.22
                 0.50 1.54 0.48 1.54 0.48 3.10 2.18 3.10 ;
    END
END latnrsqb_1

MACRO latnrsq_4
    CLASS CORE ;
    FOREIGN latnrsq_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.76 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.24 2.72 3.68 3.22 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.58 2.72 14.26 2.72 14.26 2.40 14.24 2.40 14.24 2.08
                 14.58 2.08 ;
        END
    END g
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  21.42 3.25 19.65 3.25 19.65 2.93 20.64 2.93 20.64 2.72
                 21.10 2.72 21.10 1.62 19.17 1.62 19.17 1.30 21.42 1.30 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  18.08 1.22 18.59 1.86 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.90  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.71 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.76 0.90 17.69 0.90 17.69 1.28 17.37 1.28 17.37 0.90
                 14.78 0.90 14.78 1.50 14.46 1.50 14.46 0.90 12.60 0.90
                 12.60 1.28 12.28 1.28 12.28 0.90 8.24 0.90 8.24 1.24 7.92 1.24
                 7.92 0.90 1.20 0.90 1.20 1.28 0.88 1.28 0.88 0.90 0.00 0.90
                 0.00 -0.90 21.76 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.76 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.16 1.20 4.16
                 1.20 4.86 1.56 4.86 1.56 4.16 1.88 4.16 1.88 4.86 12.28 4.86
                 12.28 4.16 12.60 4.16 12.60 4.86 14.42 4.86 14.42 4.16
                 15.30 4.16 15.30 4.86 16.67 4.86 16.67 2.95 16.99 2.95
                 16.99 4.86 20.31 4.86 20.31 4.79 20.73 4.79 20.73 4.86
                 21.76 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  18.73 2.23 19.05 3.90 ;
        POLYGON  17.75 4.54 17.43 4.54 17.43 2.52 16.21 2.52 16.21 3.84
                 15.89 3.84 15.89 2.18 15.46 2.18 15.28 2.00 15.28 1.22
                 15.60 1.22 15.60 1.86 16.21 1.86 16.21 2.20 17.75 2.20 ;
        RECT  15.98 1.22 16.99 1.54 ;
        POLYGON  15.22 3.84 5.34 3.84 5.34 4.30 5.02 4.30 5.02 3.84 4.70 3.84
                 4.70 1.90 5.02 1.90 5.02 3.52 14.90 3.52 14.90 2.40 15.22 2.40 ;
        POLYGON  14.08 1.54 13.94 1.54 13.94 1.95 13.82 2.07 13.82 2.48
                 13.94 2.60 13.94 2.88 13.98 2.88 13.98 3.20 13.62 3.20
                 13.62 2.74 13.50 2.62 13.50 1.93 13.62 1.81 13.62 1.22
                 14.08 1.22 ;
        POLYGON  13.30 1.62 13.18 1.74 13.18 2.88 13.30 2.88 13.30 3.20
                 5.34 3.20 5.34 2.44 5.66 2.44 5.66 2.88 12.86 2.88 12.86 1.47
                 12.91 1.47 12.91 1.37 12.98 1.37 12.98 1.30 13.30 1.30 ;
        POLYGON  11.92 1.60 11.60 1.60 11.60 1.54 8.88 1.54 8.88 1.88 7.28 1.88
                 7.28 1.60 6.46 1.60 6.46 1.28 7.60 1.28 7.60 1.56 8.56 1.56
                 8.56 1.22 11.92 1.22 ;
        POLYGON  11.92 4.54 5.72 4.54 5.72 4.16 6.04 4.16 6.04 4.22 11.92 4.22 ;
        POLYGON  11.22 2.52 8.70 2.52 8.70 2.20 10.90 2.20 10.90 2.04
                 11.22 2.04 ;
        POLYGON  7.46 2.52 6.46 2.52 5.82 1.88 5.82 1.54 4.38 1.54 4.38 2.24
                 2.04 2.24 2.04 1.22 2.36 1.22 2.36 1.92 4.06 1.92 4.06 1.22
                 6.14 1.22 6.14 1.74 6.60 2.20 7.46 2.20 ;
        POLYGON  4.64 4.50 3.96 4.50 3.96 4.54 3.64 4.54 3.64 4.18 4.64 4.18 ;
        POLYGON  3.74 1.60 3.42 1.60 3.42 1.54 2.74 1.54 2.74 1.22 3.74 1.22 ;
        RECT  2.26 4.22 3.26 4.54 ;
        POLYGON  2.18 3.42 0.50 3.42 0.50 4.48 0.16 4.48 0.16 1.22 0.50 1.22
                 0.50 1.54 0.48 1.54 0.48 3.10 2.18 3.10 ;
    END
END latnrsq_4

MACRO latnrsq_2
    CLASS CORE ;
    FOREIGN latnrsq_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 20.48 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.24 2.72 3.68 3.22 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.58 2.72 14.26 2.72 14.26 2.40 14.24 2.40 14.24 2.08
                 14.58 2.08 ;
        END
    END g
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.32 1.76 20.27 1.76 20.27 4.54 19.95 4.54 19.95 1.22
                 20.27 1.22 20.27 1.44 20.32 1.44 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  18.08 1.22 18.59 1.86 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.90  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.71 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 0.90 19.57 0.90 19.57 1.26 19.25 1.26 19.25 0.90
                 17.69 0.90 17.69 1.28 17.37 1.28 17.37 0.90 14.78 0.90
                 14.78 1.50 14.46 1.50 14.46 0.90 12.60 0.90 12.60 1.28
                 12.28 1.28 12.28 0.90 8.24 0.90 8.24 1.24 7.92 1.24 7.92 0.90
                 1.20 0.90 1.20 1.28 0.88 1.28 0.88 0.90 0.00 0.90 0.00 -0.90
                 20.48 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.16 1.20 4.16
                 1.20 4.86 1.56 4.86 1.56 4.16 1.88 4.16 1.88 4.86 12.28 4.86
                 12.28 4.16 12.60 4.16 12.60 4.86 14.42 4.86 14.42 4.16
                 15.30 4.16 15.30 4.86 16.67 4.86 16.67 2.95 16.99 2.95
                 16.99 4.86 19.25 4.86 19.25 4.22 19.57 4.22 19.57 4.86
                 20.48 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  19.05 3.08 18.89 3.08 18.89 4.54 18.57 4.54 18.57 2.76
                 19.05 2.76 ;
        POLYGON  17.75 4.54 17.43 4.54 17.43 2.52 16.21 2.52 16.21 3.84
                 15.89 3.84 15.89 2.18 15.46 2.18 15.28 2.00 15.28 1.22
                 15.60 1.22 15.60 1.86 16.21 1.86 16.21 2.20 17.75 2.20 ;
        RECT  15.98 1.22 16.99 1.54 ;
        POLYGON  15.22 3.84 5.34 3.84 5.34 4.30 5.02 4.30 5.02 3.84 4.70 3.84
                 4.70 1.90 5.02 1.90 5.02 3.52 14.90 3.52 14.90 2.40 15.22 2.40 ;
        POLYGON  14.08 1.54 13.94 1.54 13.94 1.95 13.82 2.07 13.82 2.48
                 13.94 2.60 13.94 2.88 13.98 2.88 13.98 3.20 13.62 3.20
                 13.62 2.74 13.50 2.62 13.50 1.93 13.62 1.81 13.62 1.22
                 14.08 1.22 ;
        POLYGON  13.30 1.62 13.18 1.74 13.18 2.88 13.30 2.88 13.30 3.20
                 5.34 3.20 5.34 2.44 5.66 2.44 5.66 2.88 12.86 2.88 12.86 1.47
                 12.91 1.47 12.91 1.37 12.98 1.37 12.98 1.30 13.30 1.30 ;
        POLYGON  11.92 1.60 11.60 1.60 11.60 1.54 8.88 1.54 8.88 1.88 7.28 1.88
                 7.28 1.60 6.46 1.60 6.46 1.28 7.60 1.28 7.60 1.56 8.56 1.56
                 8.56 1.22 11.92 1.22 ;
        POLYGON  11.92 4.54 5.72 4.54 5.72 4.16 6.04 4.16 6.04 4.22 11.92 4.22 ;
        POLYGON  11.22 2.52 8.70 2.52 8.70 2.20 10.90 2.20 10.90 2.04
                 11.22 2.04 ;
        POLYGON  7.46 2.52 6.46 2.52 5.82 1.88 5.82 1.54 4.38 1.54 4.38 2.24
                 2.04 2.24 2.04 1.22 2.36 1.22 2.36 1.92 4.06 1.92 4.06 1.22
                 6.14 1.22 6.14 1.74 6.60 2.20 7.46 2.20 ;
        POLYGON  4.64 4.50 3.96 4.50 3.96 4.54 3.64 4.54 3.64 4.18 4.64 4.18 ;
        POLYGON  3.74 1.60 3.42 1.60 3.42 1.54 2.74 1.54 2.74 1.22 3.74 1.22 ;
        RECT  2.26 4.22 3.26 4.54 ;
        POLYGON  2.18 3.42 0.50 3.42 0.50 4.48 0.16 4.48 0.16 1.22 0.50 1.22
                 0.50 1.54 0.48 1.54 0.48 3.10 2.18 3.10 ;
    END
END latnrsq_2

MACRO latnrsq_1
    CLASS CORE ;
    FOREIGN latnrsq_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 20.48 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.24 2.72 3.68 3.22 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.58 2.72 14.26 2.72 14.26 2.40 14.24 2.40 14.24 2.08
                 14.58 2.08 ;
        END
    END g
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.32 1.76 20.27 1.76 20.27 4.54 19.95 4.54 19.95 1.22
                 20.27 1.22 20.27 1.44 20.32 1.44 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  18.08 1.22 18.59 1.86 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.90  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.71 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 0.90 19.57 0.90 19.57 1.26 19.25 1.26 19.25 0.90
                 17.69 0.90 17.69 1.28 17.37 1.28 17.37 0.90 14.78 0.90
                 14.78 1.50 14.46 1.50 14.46 0.90 12.60 0.90 12.60 1.28
                 12.28 1.28 12.28 0.90 8.24 0.90 8.24 1.24 7.92 1.24 7.92 0.90
                 1.20 0.90 1.20 1.28 0.88 1.28 0.88 0.90 0.00 0.90 0.00 -0.90
                 20.48 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.16 1.20 4.16
                 1.20 4.86 1.56 4.86 1.56 4.16 1.88 4.16 1.88 4.86 12.28 4.86
                 12.28 4.16 12.60 4.16 12.60 4.86 14.42 4.86 14.42 4.16
                 15.30 4.16 15.30 4.86 16.67 4.86 16.67 2.95 16.99 2.95
                 16.99 4.86 19.25 4.86 19.25 4.22 19.57 4.22 19.57 4.86
                 20.48 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  19.05 3.08 18.89 3.08 18.89 4.54 18.57 4.54 18.57 2.76
                 19.05 2.76 ;
        POLYGON  17.75 4.54 17.43 4.54 17.43 2.52 16.21 2.52 16.21 3.84
                 15.89 3.84 15.89 2.18 15.46 2.18 15.28 2.00 15.28 1.22
                 15.60 1.22 15.60 1.86 16.21 1.86 16.21 2.20 17.75 2.20 ;
        RECT  15.98 1.22 16.99 1.54 ;
        POLYGON  15.22 3.84 5.34 3.84 5.34 4.30 5.02 4.30 5.02 3.84 4.70 3.84
                 4.70 1.90 5.02 1.90 5.02 3.52 14.90 3.52 14.90 2.40 15.22 2.40 ;
        POLYGON  14.08 1.54 13.94 1.54 13.94 1.95 13.82 2.07 13.82 2.48
                 13.94 2.60 13.94 2.88 13.98 2.88 13.98 3.20 13.62 3.20
                 13.62 2.74 13.50 2.62 13.50 1.93 13.62 1.81 13.62 1.22
                 14.08 1.22 ;
        POLYGON  13.30 1.62 13.18 1.74 13.18 2.88 13.30 2.88 13.30 3.20
                 5.34 3.20 5.34 2.44 5.66 2.44 5.66 2.88 12.86 2.88 12.86 1.47
                 12.91 1.47 12.91 1.37 12.98 1.37 12.98 1.30 13.30 1.30 ;
        POLYGON  11.92 1.60 11.60 1.60 11.60 1.54 8.88 1.54 8.88 1.88 7.28 1.88
                 7.28 1.60 6.46 1.60 6.46 1.28 7.60 1.28 7.60 1.56 8.56 1.56
                 8.56 1.22 11.92 1.22 ;
        POLYGON  11.92 4.54 5.72 4.54 5.72 4.16 6.04 4.16 6.04 4.22 11.92 4.22 ;
        POLYGON  11.22 2.52 8.70 2.52 8.70 2.20 10.90 2.20 10.90 2.04
                 11.22 2.04 ;
        POLYGON  7.46 2.52 6.46 2.52 5.82 1.88 5.82 1.54 4.38 1.54 4.38 2.24
                 2.04 2.24 2.04 1.22 2.36 1.22 2.36 1.92 4.06 1.92 4.06 1.22
                 6.14 1.22 6.14 1.74 6.60 2.20 7.46 2.20 ;
        POLYGON  4.64 4.50 3.96 4.50 3.96 4.54 3.64 4.54 3.64 4.18 4.64 4.18 ;
        POLYGON  3.74 1.60 3.42 1.60 3.42 1.54 2.74 1.54 2.74 1.22 3.74 1.22 ;
        RECT  2.26 4.22 3.26 4.54 ;
        POLYGON  2.18 3.42 0.50 3.42 0.50 4.48 0.16 4.48 0.16 1.22 0.50 1.22
                 0.50 1.54 0.48 1.54 0.48 3.10 2.18 3.10 ;
    END
END latnrsq_1

MACRO latnrs_4
    CLASS CORE ;
    FOREIGN latnrs_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.24 2.72 3.68 3.22 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.58 2.72 14.26 2.72 14.26 2.40 14.24 2.40 14.24 2.08
                 14.58 2.08 ;
        END
    END g
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  21.42 3.25 19.65 3.25 19.65 2.93 20.64 2.93 20.64 2.72
                 21.10 2.72 21.10 1.62 19.17 1.62 19.17 1.30 21.42 1.30 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  23.52 4.53 21.74 4.53 21.74 4.21 23.20 4.21 23.20 1.90
                 21.74 1.90 21.74 1.58 23.52 1.58 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  18.08 1.22 18.59 1.86 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.90  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.71 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  23.68 0.90 22.76 0.90 22.76 1.23 22.44 1.23 22.44 0.90
                 17.69 0.90 17.69 1.28 17.37 1.28 17.37 0.90 14.78 0.90
                 14.78 1.50 14.46 1.50 14.46 0.90 12.60 0.90 12.60 1.28
                 12.28 1.28 12.28 0.90 8.24 0.90 8.24 1.24 7.92 1.24 7.92 0.90
                 1.20 0.90 1.20 1.28 0.88 1.28 0.88 0.90 0.00 0.90 0.00 -0.90
                 23.68 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  23.68 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.16 1.20 4.16
                 1.20 4.86 1.56 4.86 1.56 4.16 1.88 4.16 1.88 4.86 12.28 4.86
                 12.28 4.16 12.60 4.16 12.60 4.86 14.42 4.86 14.42 4.16
                 15.30 4.16 15.30 4.86 16.67 4.86 16.67 2.95 16.99 2.95
                 16.99 4.86 20.31 4.86 20.31 4.79 20.73 4.79 20.73 4.86
                 23.68 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  22.76 3.89 19.80 3.89 19.80 4.54 17.43 4.54 17.43 2.52
                 16.21 2.52 16.21 3.84 15.89 3.84 15.89 2.18 15.46 2.18
                 15.28 2.00 15.28 1.22 15.60 1.22 15.60 1.86 16.21 1.86
                 16.21 2.20 17.75 2.20 17.75 4.22 19.48 4.22 19.48 3.57
                 22.44 3.57 22.44 2.34 22.76 2.34 ;
        RECT  18.73 2.23 19.05 3.90 ;
        RECT  15.98 1.22 16.99 1.54 ;
        POLYGON  15.22 3.84 5.34 3.84 5.34 4.30 5.02 4.30 5.02 3.84 4.70 3.84
                 4.70 1.90 5.02 1.90 5.02 3.52 14.90 3.52 14.90 2.40 15.22 2.40 ;
        POLYGON  14.08 1.54 13.94 1.54 13.94 1.95 13.82 2.07 13.82 2.48
                 13.94 2.60 13.94 2.88 13.98 2.88 13.98 3.20 13.62 3.20
                 13.62 2.74 13.50 2.62 13.50 1.93 13.62 1.81 13.62 1.22
                 14.08 1.22 ;
        POLYGON  13.30 1.62 13.18 1.74 13.18 2.88 13.30 2.88 13.30 3.20
                 5.34 3.20 5.34 2.44 5.66 2.44 5.66 2.88 12.86 2.88 12.86 1.47
                 12.91 1.47 12.91 1.37 12.98 1.37 12.98 1.30 13.30 1.30 ;
        POLYGON  11.92 1.60 11.60 1.60 11.60 1.54 8.88 1.54 8.88 1.88 7.28 1.88
                 7.28 1.60 6.46 1.60 6.46 1.28 7.60 1.28 7.60 1.56 8.56 1.56
                 8.56 1.22 11.92 1.22 ;
        POLYGON  11.92 4.54 5.72 4.54 5.72 4.16 6.04 4.16 6.04 4.22 11.92 4.22 ;
        POLYGON  11.22 2.52 8.70 2.52 8.70 2.20 10.90 2.20 10.90 2.04
                 11.22 2.04 ;
        POLYGON  7.46 2.52 6.46 2.52 5.82 1.88 5.82 1.54 4.38 1.54 4.38 2.24
                 2.04 2.24 2.04 1.22 2.36 1.22 2.36 1.92 4.06 1.92 4.06 1.22
                 6.14 1.22 6.14 1.74 6.60 2.20 7.46 2.20 ;
        POLYGON  4.64 4.50 3.96 4.50 3.96 4.54 3.64 4.54 3.64 4.18 4.64 4.18 ;
        POLYGON  3.74 1.60 3.42 1.60 3.42 1.54 2.74 1.54 2.74 1.22 3.74 1.22 ;
        RECT  2.26 4.22 3.26 4.54 ;
        POLYGON  2.18 3.42 0.50 3.42 0.50 4.48 0.16 4.48 0.16 1.22 0.50 1.22
                 0.50 1.54 0.48 1.54 0.48 3.10 2.18 3.10 ;
    END
END latnrs_4

MACRO latnrs_2
    CLASS CORE ;
    FOREIGN latnrs_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.76 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.24 2.72 3.68 3.22 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.58 2.72 14.26 2.72 14.26 2.40 14.24 2.40 14.24 2.08
                 14.58 2.08 ;
        END
    END g
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.84  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  19.73 1.76 19.69 1.76 19.69 3.37 19.73 3.37 19.73 3.69
                 19.37 3.69 19.37 1.76 19.36 1.76 19.36 1.44 19.37 1.44
                 19.37 1.22 19.73 1.22 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.71  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  21.60 2.40 21.25 2.40 21.25 3.79 20.91 3.79 20.91 3.47
                 20.93 3.47 20.93 1.54 20.81 1.54 20.81 1.22 21.25 1.22
                 21.25 2.08 21.60 2.08 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  18.08 1.22 18.59 1.86 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.90  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.71 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.76 0.90 20.43 0.90 20.43 1.36 20.11 1.36 20.11 0.90
                 17.69 0.90 17.69 1.28 17.37 1.28 17.37 0.90 14.78 0.90
                 14.78 1.14 14.46 1.14 14.46 0.90 12.60 0.90 12.60 1.28
                 12.28 1.28 12.28 0.90 8.24 0.90 8.24 1.24 7.92 1.24 7.92 0.90
                 1.20 0.90 1.20 1.58 0.88 1.58 0.88 0.90 0.00 0.90 0.00 -0.90
                 21.76 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.76 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.16 1.20 4.16
                 1.20 4.86 1.56 4.86 1.56 4.16 1.88 4.16 1.88 4.86 12.28 4.86
                 12.28 4.16 12.60 4.16 12.60 4.86 14.42 4.86 14.42 4.16
                 15.30 4.16 15.30 4.86 16.67 4.86 16.67 2.95 16.99 2.95
                 16.99 4.86 21.76 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.59 4.54 17.43 4.54 17.43 2.52 16.21 2.52 16.21 3.84
                 15.89 3.84 15.89 2.18 15.46 2.18 15.28 2.00 15.28 1.22
                 15.60 1.22 15.60 1.86 16.21 1.86 16.21 2.20 17.75 2.20
                 17.75 4.22 20.27 4.22 20.27 2.28 20.59 2.28 ;
        RECT  18.73 2.76 19.05 3.90 ;
        RECT  15.98 1.22 16.99 1.54 ;
        POLYGON  15.22 3.84 5.34 3.84 5.34 4.30 5.02 4.30 5.02 3.84 4.70 3.84
                 4.70 1.90 5.02 1.90 5.02 3.52 14.90 3.52 14.90 2.40 15.22 2.40 ;
        POLYGON  14.08 1.54 13.94 1.54 13.94 1.95 13.82 2.07 13.82 2.48
                 13.94 2.60 13.94 2.88 13.98 2.88 13.98 3.20 13.62 3.20
                 13.62 2.74 13.50 2.62 13.50 1.93 13.62 1.81 13.62 1.22
                 14.08 1.22 ;
        POLYGON  13.30 1.62 13.18 1.74 13.18 2.88 13.30 2.88 13.30 3.20
                 5.34 3.20 5.34 2.44 5.66 2.44 5.66 2.88 12.86 2.88 12.86 1.47
                 12.91 1.47 12.91 1.37 12.98 1.37 12.98 1.30 13.30 1.30 ;
        POLYGON  11.92 1.60 11.60 1.60 11.60 1.54 8.88 1.54 8.88 1.88 7.28 1.88
                 7.28 1.60 6.46 1.60 6.46 1.28 7.60 1.28 7.60 1.56 8.56 1.56
                 8.56 1.22 11.92 1.22 ;
        POLYGON  11.92 4.54 5.72 4.54 5.72 4.16 6.04 4.16 6.04 4.22 11.92 4.22 ;
        POLYGON  11.22 2.52 8.70 2.52 8.70 2.20 10.90 2.20 10.90 2.04
                 11.22 2.04 ;
        POLYGON  7.46 2.52 6.46 2.52 5.82 1.88 5.82 1.54 4.38 1.54 4.38 2.24
                 2.04 2.24 2.04 1.22 2.36 1.22 2.36 1.92 4.06 1.92 4.06 1.22
                 6.14 1.22 6.14 1.74 6.60 2.20 7.46 2.20 ;
        POLYGON  4.64 4.50 3.96 4.50 3.96 4.54 3.64 4.54 3.64 4.18 4.64 4.18 ;
        POLYGON  3.74 1.60 3.42 1.60 3.42 1.54 2.74 1.54 2.74 1.22 3.74 1.22 ;
        RECT  2.26 4.22 3.26 4.54 ;
        POLYGON  2.18 3.42 0.50 3.42 0.50 4.48 0.16 4.48 0.16 1.22 0.50 1.22
                 0.50 1.54 0.48 1.54 0.48 3.10 2.18 3.10 ;
    END
END latnrs_2

MACRO latnrs_1
    CLASS CORE ;
    FOREIGN latnrs_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.76 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.24 2.72 3.68 3.22 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.58 2.72 14.26 2.72 14.26 2.40 14.24 2.40 14.24 2.08
                 14.58 2.08 ;
        END
    END g
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.34  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  19.73 1.76 19.69 1.76 19.69 3.58 19.73 3.58 19.73 3.90
                 19.37 3.90 19.37 1.76 19.36 1.76 19.36 1.44 19.37 1.44
                 19.37 1.22 19.73 1.22 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.23  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  21.60 2.40 21.25 2.40 21.25 4.54 20.91 4.54 20.91 4.22
                 20.93 4.22 20.93 1.54 20.81 1.54 20.81 1.22 21.25 1.22
                 21.25 2.08 21.60 2.08 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  18.08 1.22 18.59 1.86 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.90  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.71 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.76 0.90 20.43 0.90 20.43 1.66 20.11 1.66 20.11 0.90
                 17.69 0.90 17.69 1.28 17.37 1.28 17.37 0.90 14.78 0.90
                 14.78 1.14 14.46 1.14 14.46 0.90 12.60 0.90 12.60 1.28
                 12.28 1.28 12.28 0.90 8.24 0.90 8.24 1.24 7.92 1.24 7.92 0.90
                 1.20 0.90 1.20 1.58 0.88 1.58 0.88 0.90 0.00 0.90 0.00 -0.90
                 21.76 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.76 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.16 1.20 4.16
                 1.20 4.86 1.56 4.86 1.56 4.16 1.88 4.16 1.88 4.86 12.28 4.86
                 12.28 4.16 12.60 4.16 12.60 4.86 14.42 4.86 14.42 4.16
                 15.30 4.16 15.30 4.86 16.67 4.86 16.67 2.95 16.99 2.95
                 16.99 4.86 21.76 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.59 4.54 17.43 4.54 17.43 2.52 16.21 2.52 16.21 3.84
                 15.89 3.84 15.89 2.18 15.46 2.18 15.28 2.00 15.28 1.22
                 15.60 1.22 15.60 1.86 16.21 1.86 16.21 2.20 17.75 2.20
                 17.75 4.22 20.27 4.22 20.27 2.28 20.59 2.28 ;
        RECT  18.73 2.76 19.05 3.90 ;
        RECT  15.98 1.22 16.99 1.54 ;
        POLYGON  15.22 3.84 5.34 3.84 5.34 4.30 5.02 4.30 5.02 3.84 4.70 3.84
                 4.70 1.90 5.02 1.90 5.02 3.52 14.90 3.52 14.90 2.40 15.22 2.40 ;
        POLYGON  14.08 1.54 13.94 1.54 13.94 1.95 13.82 2.07 13.82 2.48
                 13.94 2.60 13.94 2.88 13.98 2.88 13.98 3.20 13.62 3.20
                 13.62 2.74 13.50 2.62 13.50 1.93 13.62 1.81 13.62 1.22
                 14.08 1.22 ;
        POLYGON  13.30 1.62 13.18 1.74 13.18 2.88 13.30 2.88 13.30 3.20
                 5.34 3.20 5.34 2.44 5.66 2.44 5.66 2.88 12.86 2.88 12.86 1.47
                 12.91 1.47 12.91 1.37 12.98 1.37 12.98 1.30 13.30 1.30 ;
        POLYGON  11.92 1.60 11.60 1.60 11.60 1.54 8.88 1.54 8.88 1.88 7.28 1.88
                 7.28 1.60 6.46 1.60 6.46 1.28 7.60 1.28 7.60 1.56 8.56 1.56
                 8.56 1.22 11.92 1.22 ;
        POLYGON  11.92 4.54 5.72 4.54 5.72 4.16 6.04 4.16 6.04 4.22 11.92 4.22 ;
        POLYGON  11.22 2.52 8.70 2.52 8.70 2.20 10.90 2.20 10.90 2.04
                 11.22 2.04 ;
        POLYGON  7.46 2.52 6.46 2.52 5.82 1.88 5.82 1.54 4.38 1.54 4.38 2.24
                 2.04 2.24 2.04 1.22 2.36 1.22 2.36 1.92 4.06 1.92 4.06 1.22
                 6.14 1.22 6.14 1.74 6.60 2.20 7.46 2.20 ;
        POLYGON  4.64 4.50 3.96 4.50 3.96 4.54 3.64 4.54 3.64 4.18 4.64 4.18 ;
        POLYGON  3.74 1.60 3.42 1.60 3.42 1.54 2.74 1.54 2.74 1.22 3.74 1.22 ;
        RECT  2.26 4.22 3.26 4.54 ;
        POLYGON  2.18 3.42 0.50 3.42 0.50 4.48 0.16 4.48 0.16 1.22 0.50 1.22
                 0.50 1.54 0.48 1.54 0.48 3.10 2.18 3.10 ;
    END
END latnrs_1

MACRO latnrqb_4
    CLASS CORE ;
    FOREIGN latnrqb_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 13.44 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 4.00 2.57 4.46 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.82 3.04 ;
        END
    END g
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  13.28 4.53 11.40 4.53 11.40 4.21 12.96 4.21 12.96 1.58
                 11.40 1.58 11.40 1.26 13.28 1.26 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.94 1.94 11.38 2.58 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  13.44 0.90 10.10 0.90 10.10 1.14 9.78 1.14 9.78 0.90 1.46 0.90
                 1.46 1.42 1.14 1.42 1.14 0.90 0.00 0.90 0.00 -0.90 13.44 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  13.44 6.66 0.00 6.66 0.00 4.86 1.14 4.86 1.14 4.22 1.46 4.22
                 1.46 4.86 13.44 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  12.42 3.89 10.62 3.89 10.62 4.22 11.04 4.22 11.04 4.54
                 10.30 4.54 10.30 3.90 8.98 3.90 8.98 3.26 8.46 3.26 8.46 2.94
                 9.30 2.94 9.30 3.58 10.30 3.58 10.30 1.40 10.48 1.22
                 10.80 1.22 10.80 1.55 10.62 1.55 10.62 3.57 12.10 3.57
                 12.10 2.34 12.42 2.34 ;
        POLYGON  9.94 3.00 9.62 3.00 9.62 2.52 8.14 2.52 8.14 3.58 8.66 3.58
                 8.66 4.22 9.40 4.22 9.40 4.54 8.34 4.54 8.34 3.90 6.68 3.90
                 6.54 4.04 6.54 4.54 6.22 4.54 6.22 3.90 6.54 3.58 7.82 3.58
                 7.82 2.52 7.08 2.52 6.32 1.76 6.32 1.22 6.64 1.22 6.64 1.62
                 7.22 2.20 9.94 2.20 ;
        RECT  8.40 1.22 9.40 1.54 ;
        RECT  7.02 1.22 8.02 1.54 ;
        RECT  6.92 4.22 8.02 4.54 ;
        POLYGON  6.30 3.00 5.40 3.90 4.30 3.90 4.30 4.54 3.28 4.54 3.28 4.22
                 3.98 4.22 3.98 3.58 5.26 3.58 5.98 2.86 5.98 2.34 5.82 2.18
                 2.70 2.18 2.70 1.86 5.96 1.86 6.30 2.20 ;
        RECT  4.94 1.22 5.94 1.54 ;
        RECT  4.84 4.22 5.84 4.54 ;
        POLYGON  5.42 2.96 3.66 2.96 3.66 3.68 0.76 3.68 0.76 4.54 0.44 4.54
                 0.44 3.36 1.14 3.36 1.14 2.18 0.36 2.18 0.36 1.86 1.46 1.86
                 1.46 3.36 3.34 3.36 3.34 2.64 5.42 2.64 ;
        POLYGON  4.56 1.54 2.38 1.54 2.38 2.58 2.92 2.58 2.92 2.90 2.06 2.90
                 2.06 1.22 4.56 1.22 ;
    END
END latnrqb_4

MACRO latnrqb_2
    CLASS CORE ;
    FOREIGN latnrqb_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.80 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 4.00 2.57 4.46 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.82 3.04 ;
        END
    END g
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.88  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.64 4.54 12.22 4.54 12.22 4.22 12.32 4.22 12.32 1.75
                 12.21 1.75 12.21 1.43 12.64 1.43 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  11.04 1.94 11.36 2.58 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  12.80 0.90 10.10 0.90 10.10 1.14 9.78 1.14 9.78 0.90 1.46 0.90
                 1.46 1.42 1.14 1.42 1.14 0.90 0.00 0.90 0.00 -0.90 12.80 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  12.80 6.66 0.00 6.66 0.00 4.86 1.14 4.86 1.14 4.22 1.46 4.22
                 1.46 4.86 12.80 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  12.00 3.82 11.28 4.54 10.40 4.54 10.40 3.90 8.98 3.90
                 8.98 3.26 8.46 3.26 8.46 2.94 9.30 2.94 9.30 3.58 10.40 3.58
                 10.40 1.30 10.48 1.22 10.80 1.22 10.80 1.54 10.72 1.54
                 10.72 4.22 11.14 4.22 11.68 3.68 11.68 2.14 12.00 2.14 ;
        POLYGON  9.94 3.00 9.62 3.00 9.62 2.52 8.14 2.52 8.14 3.58 8.66 3.58
                 8.66 4.22 9.40 4.22 9.40 4.54 8.34 4.54 8.34 3.90 6.68 3.90
                 6.54 4.04 6.54 4.54 6.22 4.54 6.22 3.90 6.54 3.58 7.82 3.58
                 7.82 2.52 7.08 2.52 6.32 1.76 6.32 1.22 6.64 1.22 6.64 1.62
                 7.22 2.20 9.94 2.20 ;
        RECT  8.40 1.22 9.40 1.54 ;
        RECT  7.02 1.22 8.02 1.54 ;
        RECT  6.92 4.22 8.02 4.54 ;
        POLYGON  6.30 3.00 5.40 3.90 4.30 3.90 4.30 4.54 3.28 4.54 3.28 4.22
                 3.98 4.22 3.98 3.58 5.26 3.58 5.98 2.86 5.98 2.34 5.82 2.18
                 2.70 2.18 2.70 1.86 5.96 1.86 6.30 2.20 ;
        RECT  4.94 1.22 5.94 1.54 ;
        RECT  4.84 4.22 5.84 4.54 ;
        POLYGON  5.42 2.96 3.66 2.96 3.66 3.68 0.76 3.68 0.76 4.54 0.44 4.54
                 0.44 3.36 1.14 3.36 1.14 2.18 0.36 2.18 0.36 1.86 1.46 1.86
                 1.46 3.36 3.34 3.36 3.34 2.64 5.42 2.64 ;
        POLYGON  4.56 1.54 2.38 1.54 2.38 2.58 2.92 2.58 2.92 2.90 2.06 2.90
                 2.06 1.22 4.56 1.22 ;
    END
END latnrqb_2

MACRO latnrqb_1
    CLASS CORE ;
    FOREIGN latnrqb_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.80 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 4.00 2.57 4.46 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.82 3.04 ;
        END
    END g
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.35  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.64 4.54 12.22 4.54 12.22 4.22 12.32 4.22 12.32 1.54
                 12.21 1.54 12.21 1.22 12.64 1.22 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  11.04 1.94 11.36 2.58 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  12.80 0.90 10.10 0.90 10.10 1.14 9.78 1.14 9.78 0.90 1.46 0.90
                 1.46 1.42 1.14 1.42 1.14 0.90 0.00 0.90 0.00 -0.90 12.80 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  12.80 6.66 0.00 6.66 0.00 4.86 1.14 4.86 1.14 4.22 1.46 4.22
                 1.46 4.86 12.80 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  12.00 3.82 11.28 4.54 10.40 4.54 10.40 3.90 8.98 3.90
                 8.98 3.26 8.46 3.26 8.46 2.94 9.30 2.94 9.30 3.58 10.40 3.58
                 10.40 1.30 10.48 1.22 10.80 1.22 10.80 1.54 10.72 1.54
                 10.72 4.22 11.14 4.22 11.68 3.68 11.68 2.14 12.00 2.14 ;
        POLYGON  9.94 3.00 9.62 3.00 9.62 2.52 8.14 2.52 8.14 3.58 8.66 3.58
                 8.66 4.22 9.40 4.22 9.40 4.54 8.34 4.54 8.34 3.90 6.68 3.90
                 6.54 4.04 6.54 4.54 6.22 4.54 6.22 3.90 6.54 3.58 7.82 3.58
                 7.82 2.52 7.08 2.52 6.32 1.76 6.32 1.22 6.64 1.22 6.64 1.62
                 7.22 2.20 9.94 2.20 ;
        RECT  8.40 1.22 9.40 1.54 ;
        RECT  7.02 1.22 8.02 1.54 ;
        RECT  6.92 4.22 8.02 4.54 ;
        POLYGON  6.30 3.00 5.40 3.90 4.30 3.90 4.30 4.54 3.28 4.54 3.28 4.22
                 3.98 4.22 3.98 3.58 5.26 3.58 5.98 2.86 5.98 2.34 5.82 2.18
                 2.70 2.18 2.70 1.86 5.96 1.86 6.30 2.20 ;
        RECT  4.94 1.22 5.94 1.54 ;
        RECT  4.84 4.22 5.84 4.54 ;
        POLYGON  5.42 2.96 3.66 2.96 3.66 3.68 0.76 3.68 0.76 4.54 0.44 4.54
                 0.44 3.36 1.14 3.36 1.14 2.18 0.36 2.18 0.36 1.86 1.46 1.86
                 1.46 3.36 3.34 3.36 3.34 2.64 5.42 2.64 ;
        POLYGON  4.56 1.54 2.38 1.54 2.38 2.58 2.92 2.58 2.92 2.90 2.06 2.90
                 2.06 1.22 4.56 1.22 ;
    END
END latnrqb_1

MACRO latnrq_4
    CLASS CORE ;
    FOREIGN latnrq_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.08 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 4.00 2.57 4.46 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.82 3.04 ;
        END
    END g
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  13.65 3.25 11.88 3.25 11.88 2.93 12.96 2.93 12.96 2.72
                 13.33 2.72 13.33 1.62 11.40 1.62 11.40 1.30 13.65 1.30 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.94 1.94 11.36 2.58 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  14.08 0.90 10.10 0.90 10.10 1.14 9.78 1.14 9.78 0.90 1.46 0.90
                 1.46 1.42 1.14 1.42 1.14 0.90 0.00 0.90 0.00 -0.90 14.08 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  14.08 6.66 0.00 6.66 0.00 4.86 1.14 4.86 1.14 4.22 1.46 4.22
                 1.46 4.86 12.52 4.86 12.52 4.79 12.94 4.79 12.94 4.86
                 14.08 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  11.07 4.54 10.30 4.54 10.30 3.90 8.98 3.90 8.98 3.26 8.46 3.26
                 8.46 2.94 9.30 2.94 9.30 3.58 10.30 3.58 10.30 1.40 10.48 1.22
                 10.80 1.22 10.80 1.55 10.62 1.55 10.62 4.22 11.07 4.22 ;
        POLYGON  9.94 3.00 9.62 3.00 9.62 2.52 8.14 2.52 8.14 3.58 8.66 3.58
                 8.66 4.22 9.40 4.22 9.40 4.54 8.34 4.54 8.34 3.90 6.68 3.90
                 6.54 4.04 6.54 4.54 6.22 4.54 6.22 3.90 6.54 3.58 7.82 3.58
                 7.82 2.52 7.08 2.52 6.32 1.76 6.32 1.22 6.64 1.22 6.64 1.62
                 7.22 2.20 9.94 2.20 ;
        RECT  8.40 1.22 9.40 1.54 ;
        RECT  7.02 1.22 8.02 1.54 ;
        RECT  6.92 4.22 8.02 4.54 ;
        POLYGON  6.30 3.00 5.40 3.90 4.30 3.90 4.30 4.54 3.28 4.54 3.28 4.22
                 3.98 4.22 3.98 3.58 5.26 3.58 5.98 2.86 5.98 2.34 5.82 2.18
                 2.70 2.18 2.70 1.86 5.96 1.86 6.30 2.20 ;
        RECT  4.94 1.22 5.94 1.54 ;
        RECT  4.84 4.22 5.84 4.54 ;
        POLYGON  5.42 2.96 3.66 2.96 3.66 3.68 0.76 3.68 0.76 4.54 0.44 4.54
                 0.44 3.36 1.14 3.36 1.14 2.18 0.36 2.18 0.36 1.86 1.46 1.86
                 1.46 3.36 3.34 3.36 3.34 2.64 5.42 2.64 ;
        POLYGON  4.56 1.54 2.38 1.54 2.38 2.58 2.92 2.58 2.92 2.90 2.06 2.90
                 2.06 1.22 4.56 1.22 ;
    END
END latnrq_4

MACRO latnrq_2
    CLASS CORE ;
    FOREIGN latnrq_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.80 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 4.00 2.57 4.46 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.82 3.04 ;
        END
    END g
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.64 3.04 12.42 3.04 12.42 4.54 12.10 4.54 12.10 1.27
                 12.42 1.27 12.42 2.72 12.64 2.72 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.94 1.94 11.36 2.58 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  12.80 0.90 10.10 0.90 10.10 1.14 9.78 1.14 9.78 0.90 1.46 0.90
                 1.46 1.42 1.14 1.42 1.14 0.90 0.00 0.90 0.00 -0.90 12.80 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  12.80 6.66 0.00 6.66 0.00 4.86 1.14 4.86 1.14 4.22 1.46 4.22
                 1.46 4.86 11.40 4.86 11.40 4.22 11.72 4.22 11.72 4.86
                 12.80 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  11.04 4.54 10.30 4.54 10.30 3.90 8.98 3.90 8.98 3.26 8.46 3.26
                 8.46 2.94 9.30 2.94 9.30 3.58 10.30 3.58 10.30 1.40 10.48 1.22
                 10.80 1.22 10.80 1.54 10.62 1.54 10.62 4.22 11.04 4.22 ;
        POLYGON  9.94 3.00 9.62 3.00 9.62 2.52 8.14 2.52 8.14 3.58 8.66 3.58
                 8.66 4.22 9.40 4.22 9.40 4.54 8.34 4.54 8.34 3.90 6.68 3.90
                 6.54 4.04 6.54 4.54 6.22 4.54 6.22 3.90 6.54 3.58 7.82 3.58
                 7.82 2.52 7.08 2.52 6.32 1.76 6.32 1.22 6.64 1.22 6.64 1.62
                 7.22 2.20 9.94 2.20 ;
        RECT  8.40 1.22 9.40 1.54 ;
        RECT  7.02 1.22 8.02 1.54 ;
        RECT  6.92 4.22 8.02 4.54 ;
        POLYGON  6.30 3.00 5.40 3.90 4.30 3.90 4.30 4.54 3.28 4.54 3.28 4.22
                 3.98 4.22 3.98 3.58 5.26 3.58 5.98 2.86 5.98 2.34 5.82 2.18
                 2.70 2.18 2.70 1.86 5.96 1.86 6.30 2.20 ;
        RECT  4.94 1.22 5.94 1.54 ;
        RECT  4.84 4.22 5.84 4.54 ;
        POLYGON  5.42 2.96 3.66 2.96 3.66 3.68 0.76 3.68 0.76 4.54 0.44 4.54
                 0.44 3.36 1.14 3.36 1.14 2.18 0.36 2.18 0.36 1.86 1.46 1.86
                 1.46 3.36 3.34 3.36 3.34 2.64 5.42 2.64 ;
        POLYGON  4.56 1.54 2.38 1.54 2.38 2.58 2.92 2.58 2.92 2.90 2.06 2.90
                 2.06 1.22 4.56 1.22 ;
    END
END latnrq_2

MACRO latnrq_1
    CLASS CORE ;
    FOREIGN latnrq_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.80 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 4.00 2.57 4.46 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.82 3.04 ;
        END
    END g
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.64 3.04 12.42 3.04 12.42 4.54 12.10 4.54 12.10 1.22
                 12.42 1.22 12.42 2.72 12.64 2.72 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  11.04 1.94 11.36 2.58 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  12.80 0.90 11.72 0.90 11.72 1.54 11.40 1.54 11.40 0.90
                 10.10 0.90 10.10 1.14 9.78 1.14 9.78 0.90 1.46 0.90 1.46 1.42
                 1.14 1.42 1.14 0.90 0.00 0.90 0.00 -0.90 12.80 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  12.80 6.66 0.00 6.66 0.00 4.86 1.14 4.86 1.14 4.22 1.46 4.22
                 1.46 4.86 11.40 4.86 11.40 4.22 11.72 4.22 11.72 4.86
                 12.80 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  11.04 4.54 10.40 4.54 10.40 3.90 8.98 3.90 8.98 3.26 8.46 3.26
                 8.46 2.94 9.30 2.94 9.30 3.58 10.40 3.58 10.40 1.30 10.48 1.22
                 10.80 1.22 10.80 1.54 10.72 1.54 10.72 4.22 11.04 4.22 ;
        POLYGON  9.94 3.00 9.62 3.00 9.62 2.52 8.14 2.52 8.14 3.58 8.66 3.58
                 8.66 4.22 9.40 4.22 9.40 4.54 8.34 4.54 8.34 3.90 6.68 3.90
                 6.54 4.04 6.54 4.54 6.22 4.54 6.22 3.90 6.54 3.58 7.82 3.58
                 7.82 2.52 7.08 2.52 6.32 1.76 6.32 1.22 6.64 1.22 6.64 1.62
                 7.22 2.20 9.94 2.20 ;
        RECT  8.40 1.22 9.40 1.54 ;
        RECT  7.02 1.22 8.02 1.54 ;
        RECT  6.92 4.22 8.02 4.54 ;
        POLYGON  6.30 3.00 5.40 3.90 4.30 3.90 4.30 4.54 3.28 4.54 3.28 4.22
                 3.98 4.22 3.98 3.58 5.26 3.58 5.98 2.86 5.98 2.34 5.82 2.18
                 2.70 2.18 2.70 1.86 5.96 1.86 6.30 2.20 ;
        RECT  4.94 1.22 5.94 1.54 ;
        RECT  4.84 4.22 5.84 4.54 ;
        POLYGON  5.42 2.96 3.66 2.96 3.66 3.68 0.76 3.68 0.76 4.54 0.44 4.54
                 0.44 3.36 1.14 3.36 1.14 2.18 0.36 2.18 0.36 1.86 1.46 1.86
                 1.46 3.36 3.34 3.36 3.34 2.64 5.42 2.64 ;
        POLYGON  4.56 1.54 2.38 1.54 2.38 2.58 2.92 2.58 2.92 2.90 2.06 2.90
                 2.06 1.22 4.56 1.22 ;
    END
END latnrq_1

MACRO latnr_4
    CLASS CORE ;
    FOREIGN latnr_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.00 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 4.00 2.57 4.46 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.82 3.04 ;
        END
    END g
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  13.65 3.25 11.88 3.25 11.88 2.93 12.96 2.93 12.96 2.72
                 13.33 2.72 13.33 1.62 11.40 1.62 11.40 1.30 13.65 1.30 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  15.84 4.53 13.97 4.53 13.97 4.21 15.52 4.21 15.52 1.90
                 13.97 1.90 13.97 1.58 15.84 1.58 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.94 1.94 11.36 2.58 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 0.90 14.99 0.90 14.99 1.23 14.67 1.23 14.67 0.90
                 10.10 0.90 10.10 1.14 9.78 1.14 9.78 0.90 1.46 0.90 1.46 1.42
                 1.14 1.42 1.14 0.90 0.00 0.90 0.00 -0.90 16.00 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 6.66 0.00 6.66 0.00 4.86 1.14 4.86 1.14 4.22 1.46 4.22
                 1.46 4.86 12.52 4.86 12.52 4.79 12.94 4.79 12.94 4.86
                 16.00 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  14.99 3.89 12.64 3.89 12.64 3.90 12.00 4.54 10.30 4.54
                 10.30 3.90 8.98 3.90 8.98 3.26 8.46 3.26 8.46 2.94 9.30 2.94
                 9.30 3.58 10.30 3.58 10.30 1.40 10.48 1.22 10.80 1.22
                 10.80 1.55 10.62 1.55 10.62 4.22 11.86 4.22 12.32 3.76
                 12.32 3.57 14.67 3.57 14.67 2.34 14.99 2.34 ;
        POLYGON  9.94 3.00 9.62 3.00 9.62 2.52 8.14 2.52 8.14 3.58 8.66 3.58
                 8.66 4.22 9.40 4.22 9.40 4.54 8.34 4.54 8.34 3.90 6.68 3.90
                 6.54 4.04 6.54 4.54 6.22 4.54 6.22 3.90 6.54 3.58 7.82 3.58
                 7.82 2.52 7.08 2.52 6.32 1.76 6.32 1.22 6.64 1.22 6.64 1.62
                 7.22 2.20 9.94 2.20 ;
        RECT  8.40 1.22 9.40 1.54 ;
        RECT  7.02 1.22 8.02 1.54 ;
        RECT  6.92 4.22 8.02 4.54 ;
        POLYGON  6.30 3.00 5.40 3.90 4.30 3.90 4.30 4.54 3.28 4.54 3.28 4.22
                 3.98 4.22 3.98 3.58 5.26 3.58 5.98 2.86 5.98 2.34 5.82 2.18
                 2.70 2.18 2.70 1.86 5.96 1.86 6.30 2.20 ;
        RECT  4.94 1.22 5.94 1.54 ;
        RECT  4.84 4.22 5.84 4.54 ;
        POLYGON  5.42 2.96 3.66 2.96 3.66 3.68 0.76 3.68 0.76 4.54 0.44 4.54
                 0.44 3.36 1.14 3.36 1.14 2.18 0.36 2.18 0.36 1.86 1.46 1.86
                 1.46 3.36 3.34 3.36 3.34 2.64 5.42 2.64 ;
        POLYGON  4.56 1.54 2.38 1.54 2.38 2.58 2.92 2.58 2.92 2.90 2.06 2.90
                 2.06 1.22 4.56 1.22 ;
    END
END latnr_4

MACRO latnr_2
    CLASS CORE ;
    FOREIGN latnr_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 13.44 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 4.00 2.57 4.46 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.82 3.04 ;
        END
    END g
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.96  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.00 3.62 11.72 3.90 11.40 3.90 11.40 3.58 11.58 3.58
                 11.68 3.48 11.68 1.61 11.40 1.61 11.40 1.29 12.00 1.29 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.88  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  13.28 4.54 12.94 4.54 12.94 4.22 12.96 4.22 12.96 1.61
                 12.94 1.61 12.94 1.29 13.28 1.29 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  11.04 1.94 11.36 2.58 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  13.44 0.90 10.10 0.90 10.10 1.14 9.78 1.14 9.78 0.90 1.46 0.90
                 1.46 1.42 1.14 1.42 1.14 0.90 0.00 0.90 0.00 -0.90 13.44 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  13.44 6.66 0.00 6.66 0.00 4.86 1.14 4.86 1.14 4.22 1.46 4.22
                 1.46 4.86 13.44 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  12.64 3.90 12.00 4.54 10.40 4.54 10.40 3.90 8.98 3.90
                 8.98 3.26 8.46 3.26 8.46 2.94 9.30 2.94 9.30 3.58 10.40 3.58
                 10.40 1.30 10.48 1.22 10.80 1.22 10.80 1.54 10.72 1.54
                 10.72 4.22 11.86 4.22 12.32 3.76 12.32 2.12 12.64 2.12 ;
        POLYGON  9.94 3.00 9.62 3.00 9.62 2.52 8.14 2.52 8.14 3.58 8.66 3.58
                 8.66 4.22 9.40 4.22 9.40 4.54 8.34 4.54 8.34 3.90 6.68 3.90
                 6.54 4.04 6.54 4.54 6.22 4.54 6.22 3.90 6.54 3.58 7.82 3.58
                 7.82 2.52 7.08 2.52 6.32 1.76 6.32 1.22 6.64 1.22 6.64 1.62
                 7.22 2.20 9.94 2.20 ;
        RECT  8.40 1.22 9.40 1.54 ;
        RECT  7.02 1.22 8.02 1.54 ;
        RECT  6.92 4.22 8.02 4.54 ;
        POLYGON  6.30 3.00 5.40 3.90 4.30 3.90 4.30 4.54 3.28 4.54 3.28 4.22
                 3.98 4.22 3.98 3.58 5.26 3.58 5.98 2.86 5.98 2.34 5.82 2.18
                 2.70 2.18 2.70 1.86 5.96 1.86 6.30 2.20 ;
        RECT  4.94 1.22 5.94 1.54 ;
        RECT  4.84 4.22 5.84 4.54 ;
        POLYGON  5.42 2.96 3.66 2.96 3.66 3.68 0.76 3.68 0.76 4.54 0.44 4.54
                 0.44 3.36 1.14 3.36 1.14 2.18 0.36 2.18 0.36 1.86 1.46 1.86
                 1.46 3.36 3.34 3.36 3.34 2.64 5.42 2.64 ;
        POLYGON  4.56 1.54 2.38 1.54 2.38 2.58 2.92 2.58 2.92 2.90 2.06 2.90
                 2.06 1.22 4.56 1.22 ;
    END
END latnr_2

MACRO latnr_1
    CLASS CORE ;
    FOREIGN latnr_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 13.44 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 4.00 2.57 4.46 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.82 3.04 ;
        END
    END g
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.44  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.00 3.62 11.72 3.90 11.40 3.90 11.40 3.58 11.58 3.58
                 11.68 3.48 11.68 1.54 11.40 1.54 11.40 1.22 12.00 1.22 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.35  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  13.28 4.54 12.94 4.54 12.94 4.22 12.96 4.22 12.96 1.54
                 12.94 1.54 12.94 1.22 13.28 1.22 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  11.04 1.94 11.36 2.58 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  13.44 0.90 10.10 0.90 10.10 1.14 9.78 1.14 9.78 0.90 1.46 0.90
                 1.46 1.42 1.14 1.42 1.14 0.90 0.00 0.90 0.00 -0.90 13.44 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  13.44 6.66 0.00 6.66 0.00 4.86 1.14 4.86 1.14 4.22 1.46 4.22
                 1.46 4.86 13.44 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  12.64 3.90 12.00 4.54 10.40 4.54 10.40 3.90 8.98 3.90
                 8.98 3.26 8.46 3.26 8.46 2.94 9.30 2.94 9.30 3.58 10.40 3.58
                 10.40 1.30 10.48 1.22 10.80 1.22 10.80 1.54 10.72 1.54
                 10.72 4.22 11.86 4.22 12.32 3.76 12.32 2.14 12.64 2.14 ;
        POLYGON  9.94 3.00 9.62 3.00 9.62 2.52 8.14 2.52 8.14 3.58 8.66 3.58
                 8.66 4.22 9.40 4.22 9.40 4.54 8.34 4.54 8.34 3.90 6.68 3.90
                 6.54 4.04 6.54 4.54 6.22 4.54 6.22 3.90 6.54 3.58 7.82 3.58
                 7.82 2.52 7.08 2.52 6.32 1.76 6.32 1.22 6.64 1.22 6.64 1.62
                 7.22 2.20 9.94 2.20 ;
        RECT  8.40 1.22 9.40 1.54 ;
        RECT  7.02 1.22 8.02 1.54 ;
        RECT  6.92 4.22 8.02 4.54 ;
        POLYGON  6.30 3.00 5.40 3.90 4.30 3.90 4.30 4.54 3.28 4.54 3.28 4.22
                 3.98 4.22 3.98 3.58 5.26 3.58 5.98 2.86 5.98 2.34 5.82 2.18
                 2.70 2.18 2.70 1.86 5.96 1.86 6.30 2.20 ;
        RECT  4.94 1.22 5.94 1.54 ;
        RECT  4.84 4.22 5.84 4.54 ;
        POLYGON  5.42 2.96 3.66 2.96 3.66 3.68 0.76 3.68 0.76 4.54 0.44 4.54
                 0.44 3.36 1.14 3.36 1.14 2.18 0.36 2.18 0.36 1.86 1.46 1.86
                 1.46 3.36 3.34 3.36 3.34 2.64 5.42 2.64 ;
        POLYGON  4.56 1.54 2.38 1.54 2.38 2.58 2.92 2.58 2.92 2.90 2.06 2.90
                 2.06 1.22 4.56 1.22 ;
    END
END latnr_1

MACRO latnqb_4
    CLASS CORE ;
    FOREIGN latnqb_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.24 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.08 7.16 2.54 ;
        END
    END g
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.08 4.53 8.32 4.53 8.32 4.21 9.76 4.21 9.76 1.90 8.32 1.90
                 8.32 1.58 10.08 1.58 ;
        END
    END qb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  10.24 0.90 9.34 0.90 9.34 1.23 9.02 1.23 9.02 0.90 7.06 0.90
                 7.06 1.12 6.74 1.12 6.74 0.90 4.88 0.90 4.88 1.14 4.56 1.14
                 4.56 0.90 1.20 0.90 1.20 1.62 0.88 1.62 0.88 0.90 0.00 0.90
                 0.00 -0.90 10.24 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  10.24 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 4.66 4.86 4.66 4.62 4.98 4.62 4.98 4.86 6.74 4.86
                 6.74 4.62 7.06 4.62 7.06 4.86 10.24 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  9.34 3.89 7.76 3.89 7.76 4.45 7.44 4.45 7.44 3.42 7.54 3.42
                 7.54 1.54 7.44 1.54 7.44 1.22 7.86 1.22 7.86 3.57 9.02 3.57
                 9.02 2.30 9.34 2.30 ;
        POLYGON  7.22 3.18 7.00 3.18 7.00 4.30 4.66 4.30 4.66 3.90 2.74 3.90
                 2.74 4.54 2.42 4.54 2.42 1.30 2.74 1.30 2.74 3.58 4.98 3.58
                 4.98 3.98 6.68 3.98 6.68 2.86 7.22 2.86 ;
        POLYGON  6.36 1.54 6.32 1.54 6.32 1.80 5.97 2.15 5.97 2.71 6.32 3.06
                 6.32 3.34 6.36 3.34 6.36 3.66 6.00 3.66 6.00 3.20 5.65 2.85
                 5.65 2.01 6.00 1.66 6.00 1.22 6.36 1.22 ;
        POLYGON  5.68 3.66 5.36 3.66 5.36 3.48 5.14 3.26 4.66 3.26 4.66 3.18
                 3.06 3.18 3.06 2.86 4.66 2.86 4.66 1.90 5.26 1.30 5.58 1.30
                 5.58 1.62 5.40 1.62 4.98 2.04 4.98 2.94 5.28 2.94 5.68 3.34 ;
        RECT  3.18 4.22 4.28 4.54 ;
        RECT  3.18 1.58 4.18 1.90 ;
        POLYGON  2.00 2.26 0.18 2.26 0.18 1.30 0.50 1.30 0.50 1.94 1.68 1.94
                 1.68 1.30 2.00 1.30 ;
        POLYGON  1.88 4.54 1.56 4.54 1.56 3.76 0.50 3.76 0.50 4.54 0.18 4.54
                 0.18 3.44 1.88 3.44 ;
    END
END latnqb_4

MACRO latnqb_2
    CLASS CORE ;
    FOREIGN latnqb_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.24 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.08 7.16 2.54 ;
        END
    END g
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.08 3.72 9.46 3.72 9.46 4.38 9.14 4.38 9.14 3.40 9.76 3.40
                 9.76 1.92 9.14 1.92 9.14 1.60 10.08 1.60 ;
        END
    END qb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  10.24 0.90 8.76 0.90 8.76 1.08 8.44 1.08 8.44 0.90 7.06 0.90
                 7.06 1.12 6.74 1.12 6.74 0.90 4.88 0.90 4.88 1.14 4.56 1.14
                 4.56 0.90 1.20 0.90 1.20 1.62 0.88 1.62 0.88 0.90 0.00 0.90
                 0.00 -0.90 10.24 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  10.24 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 4.66 4.86 4.66 4.62 4.98 4.62 4.98 4.86 6.74 4.86
                 6.74 4.62 7.06 4.62 7.06 4.86 10.24 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  8.92 2.62 8.82 2.62 8.82 4.10 8.12 4.10 8.12 4.54 7.80 4.54
                 7.80 4.10 7.54 4.10 7.54 3.74 7.44 3.74 7.44 3.42 7.54 3.42
                 7.54 1.54 7.44 1.54 7.44 1.22 7.86 1.22 7.86 3.78 8.50 3.78
                 8.50 2.30 8.92 2.30 ;
        POLYGON  7.22 3.18 7.00 3.18 7.00 4.30 4.66 4.30 4.66 3.90 2.74 3.90
                 2.74 4.54 2.42 4.54 2.42 1.30 2.74 1.30 2.74 3.58 4.98 3.58
                 4.98 3.98 6.68 3.98 6.68 2.86 7.22 2.86 ;
        POLYGON  6.36 1.54 6.32 1.54 6.32 1.80 5.97 2.15 5.97 2.71 6.32 3.06
                 6.32 3.34 6.36 3.34 6.36 3.66 6.00 3.66 6.00 3.20 5.65 2.85
                 5.65 2.01 6.00 1.66 6.00 1.22 6.36 1.22 ;
        POLYGON  5.68 3.66 5.36 3.66 5.36 3.48 5.14 3.26 4.66 3.26 4.66 3.18
                 3.06 3.18 3.06 2.86 4.66 2.86 4.66 1.90 5.26 1.30 5.58 1.30
                 5.58 1.62 5.40 1.62 4.98 2.04 4.98 2.94 5.28 2.94 5.68 3.34 ;
        RECT  3.18 4.22 4.28 4.54 ;
        RECT  3.18 1.58 4.18 1.90 ;
        POLYGON  2.00 2.26 0.18 2.26 0.18 1.30 0.50 1.30 0.50 1.94 1.68 1.94
                 1.68 1.30 2.00 1.30 ;
        POLYGON  1.88 4.54 1.56 4.54 1.56 3.76 0.50 3.76 0.50 4.54 0.18 4.54
                 0.18 3.44 1.88 3.44 ;
    END
END latnqb_2

MACRO latnqb_1
    CLASS CORE ;
    FOREIGN latnqb_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.24 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.08 7.16 2.54 ;
        END
    END g
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.08 4.54 9.14 4.54 9.14 4.22 9.76 4.22 9.76 1.54 9.14 1.54
                 9.14 1.22 10.08 1.22 ;
        END
    END qb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  10.24 0.90 8.76 0.90 8.76 1.08 8.44 1.08 8.44 0.90 7.06 0.90
                 7.06 1.12 6.74 1.12 6.74 0.90 4.88 0.90 4.88 1.14 4.56 1.14
                 4.56 0.90 1.20 0.90 1.20 1.62 0.88 1.62 0.88 0.90 0.00 0.90
                 0.00 -0.90 10.24 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  10.24 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 4.66 4.86 4.66 4.62 4.98 4.62 4.98 4.86 6.74 4.86
                 6.74 4.62 7.06 4.62 7.06 4.86 8.44 4.86 8.44 4.42 8.76 4.42
                 8.76 4.86 10.24 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  8.92 2.62 8.82 2.62 8.82 4.10 8.12 4.10 8.12 4.54 7.80 4.54
                 7.80 4.10 7.54 4.10 7.54 3.74 7.44 3.74 7.44 3.42 7.54 3.42
                 7.54 1.54 7.44 1.54 7.44 1.22 7.86 1.22 7.86 3.78 8.50 3.78
                 8.50 2.30 8.92 2.30 ;
        POLYGON  7.22 3.18 7.00 3.18 7.00 4.30 4.66 4.30 4.66 3.90 2.74 3.90
                 2.74 4.54 2.42 4.54 2.42 1.30 2.74 1.30 2.74 3.58 4.98 3.58
                 4.98 3.98 6.68 3.98 6.68 2.86 7.22 2.86 ;
        POLYGON  6.36 1.54 6.32 1.54 6.32 1.80 5.97 2.15 5.97 2.71 6.32 3.06
                 6.32 3.34 6.36 3.34 6.36 3.66 6.00 3.66 6.00 3.20 5.65 2.85
                 5.65 2.01 6.00 1.66 6.00 1.22 6.36 1.22 ;
        POLYGON  5.68 3.66 5.36 3.66 5.36 3.48 5.14 3.26 4.66 3.26 4.66 3.18
                 3.06 3.18 3.06 2.86 4.66 2.86 4.66 1.90 5.26 1.30 5.58 1.30
                 5.58 1.62 5.40 1.62 4.98 2.04 4.98 2.94 5.28 2.94 5.68 3.34 ;
        RECT  3.18 4.22 4.28 4.54 ;
        RECT  3.18 1.58 4.18 1.90 ;
        POLYGON  2.00 2.26 0.18 2.26 0.18 1.30 0.50 1.30 0.50 1.94 1.68 1.94
                 1.68 1.30 2.00 1.30 ;
        POLYGON  1.88 4.54 1.56 4.54 1.56 3.76 0.50 3.76 0.50 4.54 0.18 4.54
                 0.18 3.44 1.88 3.44 ;
    END
END latnqb_1

MACRO latnq_4
    CLASS CORE ;
    FOREIGN latnq_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.24 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.08 7.16 2.54 ;
        END
    END g
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.08 3.25 8.23 3.25 8.23 2.93 9.76 2.93 9.76 1.96 8.12 1.96
                 8.12 1.64 10.08 1.64 ;
        END
    END q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  10.24 0.90 9.14 0.90 9.14 1.23 8.82 1.23 8.82 0.90 7.06 0.90
                 7.06 1.12 6.74 1.12 6.74 0.90 4.88 0.90 4.88 1.14 4.56 1.14
                 4.56 0.90 1.20 0.90 1.20 1.62 0.88 1.62 0.88 0.90 0.00 0.90
                 0.00 -0.90 10.24 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  10.24 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 4.66 4.86 4.66 4.62 4.98 4.62 4.98 4.86 6.74 4.86
                 6.74 4.62 7.06 4.62 7.06 4.86 8.87 4.86 8.87 4.79 9.29 4.79
                 9.29 4.86 10.24 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  8.12 4.54 7.80 4.54 7.80 3.89 7.44 3.89 7.44 3.42 7.54 3.42
                 7.54 2.65 7.48 2.65 7.48 1.54 7.44 1.54 7.44 1.22 7.80 1.22
                 7.80 2.33 7.86 2.33 7.86 3.57 8.12 3.57 ;
        POLYGON  7.22 3.18 7.00 3.18 7.00 4.30 4.66 4.30 4.66 3.90 2.74 3.90
                 2.74 4.54 2.42 4.54 2.42 1.30 2.74 1.30 2.74 3.58 4.98 3.58
                 4.98 3.98 6.68 3.98 6.68 2.86 7.22 2.86 ;
        POLYGON  6.36 1.54 6.32 1.54 6.32 1.80 5.97 2.15 5.97 2.71 6.32 3.06
                 6.32 3.34 6.36 3.34 6.36 3.66 6.00 3.66 6.00 3.20 5.65 2.85
                 5.65 2.01 6.00 1.66 6.00 1.22 6.36 1.22 ;
        POLYGON  5.68 3.66 5.36 3.66 5.36 3.48 5.14 3.26 4.66 3.26 4.66 3.18
                 3.06 3.18 3.06 2.86 4.66 2.86 4.66 1.90 5.26 1.30 5.58 1.30
                 5.58 1.62 5.40 1.62 4.98 2.04 4.98 2.94 5.28 2.94 5.68 3.34 ;
        RECT  3.18 4.22 4.28 4.54 ;
        RECT  3.18 1.58 4.18 1.90 ;
        POLYGON  2.00 2.26 0.18 2.26 0.18 1.30 0.50 1.30 0.50 1.94 1.68 1.94
                 1.68 1.30 2.00 1.30 ;
        POLYGON  1.88 4.54 1.56 4.54 1.56 3.76 0.50 3.76 0.50 4.54 0.18 4.54
                 0.18 3.44 1.88 3.44 ;
    END
END latnq_4

MACRO latnq_2
    CLASS CORE ;
    FOREIGN latnq_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.60 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.08 7.16 2.54 ;
        END
    END g
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.44 2.40 9.26 2.40 9.26 3.90 8.94 3.90 8.94 1.64 9.26 1.64
                 9.26 2.08 9.44 2.08 ;
        END
    END q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  9.60 0.90 8.56 0.90 8.56 1.96 8.24 1.96 8.24 0.90 7.06 0.90
                 7.06 1.12 6.74 1.12 6.74 0.90 4.88 0.90 4.88 1.14 4.56 1.14
                 4.56 0.90 1.20 0.90 1.20 1.62 0.88 1.62 0.88 0.90 0.00 0.90
                 0.00 -0.90 9.60 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  9.60 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 4.66 4.86 4.66 4.62 4.98 4.62 4.98 4.86 6.74 4.86
                 6.74 4.62 7.06 4.62 7.06 4.86 9.60 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  8.12 4.54 7.80 4.54 7.80 4.10 7.54 4.10 7.54 3.74 7.44 3.74
                 7.44 3.42 7.54 3.42 7.54 1.54 7.44 1.54 7.44 1.22 7.86 1.22
                 7.86 3.78 8.12 3.78 ;
        POLYGON  7.22 3.18 7.00 3.18 7.00 4.30 4.66 4.30 4.66 3.90 2.74 3.90
                 2.74 4.54 2.42 4.54 2.42 1.30 2.74 1.30 2.74 3.58 4.98 3.58
                 4.98 3.98 6.68 3.98 6.68 2.86 7.22 2.86 ;
        POLYGON  6.36 1.54 6.32 1.54 6.32 1.80 5.97 2.15 5.97 2.71 6.32 3.06
                 6.32 3.34 6.36 3.34 6.36 3.66 6.00 3.66 6.00 3.20 5.65 2.85
                 5.65 2.01 6.00 1.66 6.00 1.22 6.36 1.22 ;
        POLYGON  5.68 3.66 5.36 3.66 5.36 3.48 5.14 3.26 4.66 3.26 4.66 3.18
                 3.06 3.18 3.06 2.86 4.66 2.86 4.66 1.90 5.26 1.30 5.58 1.30
                 5.58 1.62 5.40 1.62 4.98 2.04 4.98 2.94 5.28 2.94 5.68 3.34 ;
        RECT  3.18 4.22 4.28 4.54 ;
        RECT  3.18 1.58 4.18 1.90 ;
        POLYGON  2.00 2.26 0.18 2.26 0.18 1.30 0.50 1.30 0.50 1.94 1.68 1.94
                 1.68 1.30 2.00 1.30 ;
        POLYGON  1.88 4.54 1.56 4.54 1.56 3.76 0.50 3.76 0.50 4.54 0.18 4.54
                 0.18 3.44 1.88 3.44 ;
    END
END latnq_2

MACRO latnq_1
    CLASS CORE ;
    FOREIGN latnq_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.60 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.08 7.16 2.54 ;
        END
    END g
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.44 2.40 9.26 2.40 9.26 4.30 8.94 4.30 8.94 1.22 9.26 1.22
                 9.26 2.08 9.44 2.08 ;
        END
    END q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  9.60 0.90 8.56 0.90 8.56 1.54 8.24 1.54 8.24 0.90 7.06 0.90
                 7.06 1.12 6.74 1.12 6.74 0.90 4.88 0.90 4.88 1.14 4.56 1.14
                 4.56 0.90 1.20 0.90 1.20 1.62 0.88 1.62 0.88 0.90 0.00 0.90
                 0.00 -0.90 9.60 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  9.60 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 4.66 4.86 4.66 4.62 4.98 4.62 4.98 4.86 6.74 4.86
                 6.74 4.62 7.06 4.62 7.06 4.86 9.60 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  8.12 4.54 7.80 4.54 7.80 4.10 7.54 4.10 7.54 3.74 7.44 3.74
                 7.44 3.42 7.54 3.42 7.54 1.54 7.44 1.54 7.44 1.22 7.86 1.22
                 7.86 3.78 8.12 3.78 ;
        POLYGON  7.22 3.18 7.00 3.18 7.00 4.30 4.66 4.30 4.66 3.90 2.74 3.90
                 2.74 4.54 2.42 4.54 2.42 1.30 2.74 1.30 2.74 3.58 4.98 3.58
                 4.98 3.98 6.68 3.98 6.68 2.86 7.22 2.86 ;
        POLYGON  6.36 1.54 6.32 1.54 6.32 1.80 5.97 2.15 5.97 2.71 6.32 3.06
                 6.32 3.34 6.36 3.34 6.36 3.66 6.00 3.66 6.00 3.20 5.65 2.85
                 5.65 2.01 6.00 1.66 6.00 1.22 6.36 1.22 ;
        POLYGON  5.68 3.66 5.36 3.66 5.36 3.48 5.14 3.26 4.66 3.26 4.66 3.18
                 3.06 3.18 3.06 2.86 4.66 2.86 4.66 1.90 5.26 1.30 5.58 1.30
                 5.58 1.62 5.40 1.62 4.98 2.04 4.98 2.94 5.28 2.94 5.68 3.34 ;
        RECT  3.18 4.22 4.28 4.54 ;
        RECT  3.18 1.58 4.18 1.90 ;
        POLYGON  2.00 2.26 0.18 2.26 0.18 1.30 0.50 1.30 0.50 1.94 1.68 1.94
                 1.68 1.30 2.00 1.30 ;
        POLYGON  1.88 4.54 1.56 4.54 1.56 3.76 0.50 3.76 0.50 4.54 0.18 4.54
                 0.18 3.44 1.88 3.44 ;
    END
END latnq_1

MACRO latn_4
    CLASS CORE ;
    FOREIGN latn_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.80 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.08 7.16 2.54 ;
        END
    END g
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.08 3.25 8.23 3.25 8.23 2.93 9.63 2.93 9.63 1.96 8.24 1.96
                 8.24 1.64 10.00 1.64 10.00 2.72 10.08 2.72 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.04 4.53 10.32 4.53 10.32 4.21 11.68 4.21 11.68 1.90
                 10.32 1.90 10.32 1.58 12.04 1.58 ;
        END
    END qb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  12.80 0.90 11.34 0.90 11.34 1.23 11.02 1.23 11.02 0.90
                 9.26 0.90 9.26 1.23 8.94 1.23 8.94 0.90 7.06 0.90 7.06 1.12
                 6.74 1.12 6.74 0.90 4.88 0.90 4.88 1.14 4.56 1.14 4.56 0.90
                 1.20 0.90 1.20 1.62 0.88 1.62 0.88 0.90 0.00 0.90 0.00 -0.90
                 12.80 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  12.80 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 4.66 4.86 4.66 4.62 4.98 4.62 4.98 4.86 6.74 4.86
                 6.74 4.62 7.06 4.62 7.06 4.86 8.87 4.86 8.87 4.79 9.29 4.79
                 9.29 4.86 12.80 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  11.34 3.89 8.12 3.89 8.12 4.54 7.80 4.54 7.80 3.89 7.54 3.89
                 7.54 3.74 7.44 3.74 7.44 3.42 7.54 3.42 7.54 1.54 7.44 1.54
                 7.44 1.22 7.86 1.22 7.86 3.57 11.02 3.57 11.02 2.30 11.34 2.30 ;
        POLYGON  7.22 3.18 7.00 3.18 7.00 4.30 4.66 4.30 4.66 3.90 2.74 3.90
                 2.74 4.54 2.42 4.54 2.42 1.30 2.74 1.30 2.74 3.58 4.98 3.58
                 4.98 3.98 6.68 3.98 6.68 2.86 7.22 2.86 ;
        POLYGON  6.36 1.54 6.32 1.54 6.32 1.80 5.97 2.15 5.97 2.71 6.32 3.06
                 6.32 3.34 6.36 3.34 6.36 3.66 6.00 3.66 6.00 3.20 5.65 2.85
                 5.65 2.01 6.00 1.66 6.00 1.22 6.36 1.22 ;
        POLYGON  5.68 3.66 5.36 3.66 5.36 3.48 5.14 3.26 4.66 3.26 4.66 3.18
                 3.06 3.18 3.06 2.86 4.66 2.86 4.66 1.90 5.26 1.30 5.58 1.30
                 5.58 1.62 5.40 1.62 4.98 2.04 4.98 2.94 5.28 2.94 5.68 3.34 ;
        RECT  3.18 4.22 4.28 4.54 ;
        RECT  3.18 1.58 4.18 1.90 ;
        POLYGON  2.00 2.26 0.18 2.26 0.18 1.30 0.50 1.30 0.50 1.94 1.68 1.94
                 1.68 1.30 2.00 1.30 ;
        POLYGON  1.88 4.54 1.56 4.54 1.56 3.76 0.50 3.76 0.50 4.54 0.18 4.54
                 0.18 3.44 1.88 3.44 ;
    END
END latn_4

MACRO latn_2
    CLASS CORE ;
    FOREIGN latn_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.24 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.08 7.16 2.54 ;
        END
    END g
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.77  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.80 1.76 8.50 1.76 8.50 3.46 8.18 3.46 8.18 1.44 8.80 1.44 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.08 3.75 9.66 3.75 9.66 3.43 9.76 3.43 9.76 1.96 9.66 1.96
                 9.66 1.64 10.08 1.64 ;
        END
    END qb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  10.24 0.90 9.28 0.90 9.28 1.08 8.96 1.08 8.96 0.90 7.06 0.90
                 7.06 1.12 6.74 1.12 6.74 0.90 4.88 0.90 4.88 1.14 4.56 1.14
                 4.56 0.90 1.20 0.90 1.20 1.62 0.88 1.62 0.88 0.90 0.00 0.90
                 0.00 -0.90 10.24 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  10.24 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 4.66 4.86 4.66 4.62 4.98 4.62 4.98 4.86 6.74 4.86
                 6.74 4.62 7.06 4.62 7.06 4.86 10.24 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  9.44 2.62 9.34 2.62 9.34 4.10 8.12 4.10 8.12 4.54 7.80 4.54
                 7.80 4.10 7.54 4.10 7.54 3.74 7.44 3.74 7.44 3.42 7.54 3.42
                 7.54 1.54 7.44 1.54 7.44 1.22 7.86 1.22 7.86 3.78 9.02 3.78
                 9.02 2.30 9.44 2.30 ;
        POLYGON  7.22 3.18 7.00 3.18 7.00 4.30 4.66 4.30 4.66 3.90 2.74 3.90
                 2.74 4.54 2.42 4.54 2.42 1.30 2.74 1.30 2.74 3.58 4.98 3.58
                 4.98 3.98 6.68 3.98 6.68 2.86 7.22 2.86 ;
        POLYGON  6.36 1.54 6.32 1.54 6.32 1.80 5.97 2.15 5.97 2.71 6.32 3.06
                 6.32 3.34 6.36 3.34 6.36 3.66 6.00 3.66 6.00 3.20 5.65 2.85
                 5.65 2.01 6.00 1.66 6.00 1.22 6.36 1.22 ;
        POLYGON  5.68 3.66 5.36 3.66 5.36 3.48 5.14 3.26 4.66 3.26 4.66 3.18
                 3.06 3.18 3.06 2.86 4.66 2.86 4.66 1.90 5.26 1.30 5.58 1.30
                 5.58 1.62 5.40 1.62 4.98 2.04 4.98 2.94 5.28 2.94 5.68 3.34 ;
        RECT  3.18 4.22 4.28 4.54 ;
        RECT  3.18 1.58 4.18 1.90 ;
        POLYGON  2.00 2.26 0.18 2.26 0.18 1.30 0.50 1.30 0.50 1.94 1.68 1.94
                 1.68 1.30 2.00 1.30 ;
        POLYGON  1.88 4.54 1.56 4.54 1.56 3.76 0.50 3.76 0.50 4.54 0.18 4.54
                 0.18 3.44 1.88 3.44 ;
    END
END latn_2

MACRO latn_1
    CLASS CORE ;
    FOREIGN latn_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.24 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END d
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.08 7.16 2.54 ;
        END
    END g
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.30  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.80 1.76 8.50 1.76 8.50 3.46 8.18 3.46 8.18 1.22 8.58 1.22
                 8.58 1.44 8.80 1.44 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.08 4.54 9.66 4.54 9.66 4.22 9.76 4.22 9.76 1.54 9.66 1.54
                 9.66 1.22 10.08 1.22 ;
        END
    END qb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  10.24 0.90 9.28 0.90 9.28 1.08 8.96 1.08 8.96 0.90 7.06 0.90
                 7.06 1.12 6.74 1.12 6.74 0.90 4.88 0.90 4.88 1.14 4.56 1.14
                 4.56 0.90 1.20 0.90 1.20 1.62 0.88 1.62 0.88 0.90 0.00 0.90
                 0.00 -0.90 10.24 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  10.24 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 4.66 4.86 4.66 4.62 4.98 4.62 4.98 4.86 6.74 4.86
                 6.74 4.62 7.06 4.62 7.06 4.86 8.96 4.86 8.96 4.42 9.28 4.42
                 9.28 4.86 10.24 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  9.44 2.62 9.34 2.62 9.34 4.10 8.12 4.10 8.12 4.54 7.80 4.54
                 7.80 4.10 7.54 4.10 7.54 3.74 7.44 3.74 7.44 3.42 7.54 3.42
                 7.54 1.54 7.44 1.54 7.44 1.22 7.86 1.22 7.86 3.78 9.02 3.78
                 9.02 2.30 9.44 2.30 ;
        POLYGON  7.22 3.18 7.00 3.18 7.00 4.30 4.66 4.30 4.66 3.90 2.74 3.90
                 2.74 4.54 2.42 4.54 2.42 1.30 2.74 1.30 2.74 3.58 4.98 3.58
                 4.98 3.98 6.68 3.98 6.68 2.86 7.22 2.86 ;
        POLYGON  6.36 1.54 6.32 1.54 6.32 1.80 5.97 2.15 5.97 2.71 6.32 3.06
                 6.32 3.34 6.36 3.34 6.36 3.66 6.00 3.66 6.00 3.20 5.65 2.85
                 5.65 2.01 6.00 1.66 6.00 1.22 6.36 1.22 ;
        POLYGON  5.68 3.66 5.36 3.66 5.36 3.48 5.14 3.26 4.66 3.26 4.66 3.18
                 3.06 3.18 3.06 2.86 4.66 2.86 4.66 1.90 5.26 1.30 5.58 1.30
                 5.58 1.62 5.40 1.62 4.98 2.04 4.98 2.94 5.28 2.94 5.68 3.34 ;
        RECT  3.18 4.22 4.28 4.54 ;
        RECT  3.18 1.58 4.18 1.90 ;
        POLYGON  2.00 2.26 0.18 2.26 0.18 1.30 0.50 1.30 0.50 1.94 1.68 1.94
                 1.68 1.30 2.00 1.30 ;
        POLYGON  1.88 4.54 1.56 4.54 1.56 3.76 0.50 3.76 0.50 4.54 0.18 4.54
                 0.18 3.44 1.88 3.44 ;
    END
END latn_1

MACRO inv_8
    CLASS CORE ;
    FOREIGN inv_8 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.84 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.72  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.34 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.29  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.30 1.96 1.90 1.96 1.90 3.78 2.98 3.78 2.98 3.10 3.30 3.10
                 3.30 4.10 0.18 4.10 0.18 3.16 0.50 3.16 0.50 3.78 1.58 3.78
                 1.58 3.04 1.44 3.04 1.44 2.72 1.58 2.72 1.58 1.96 0.18 1.96
                 0.18 1.64 3.30 1.64 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  3.84 0.90 2.60 0.90 2.60 1.32 2.28 1.32 2.28 0.90 1.20 0.90
                 1.20 1.32 0.88 1.32 0.88 0.90 0.00 0.90 0.00 -0.90 3.84 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  3.84 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.42 1.20 4.42
                 1.20 4.86 2.28 4.86 2.28 4.42 2.60 4.42 2.60 4.86 3.84 4.86 ;
        END
    END vdd!
END inv_8

MACRO inv_64
    CLASS CORE ;
    FOREIGN inv_64 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 21.77  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.34 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 32.81  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  22.90 1.96 21.50 1.96 21.50 2.72 21.60 2.72 21.60 3.04
                 21.50 3.04 21.50 3.78 22.58 3.78 22.58 3.16 22.90 3.16
                 22.90 4.10 21.18 4.10 21.18 1.96 18.70 1.96 18.70 3.78
                 19.78 3.78 19.78 3.10 20.10 3.10 20.10 3.78 21.18 3.78
                 21.18 4.10 18.38 4.10 18.38 1.96 15.90 1.96 15.90 3.78
                 16.98 3.78 16.98 3.16 17.30 3.16 17.30 3.78 18.38 3.78
                 18.38 4.10 15.58 4.10 15.58 1.96 13.10 1.96 13.10 2.72
                 13.32 2.72 13.32 3.04 13.10 3.04 13.10 3.78 14.18 3.78
                 14.18 3.10 14.50 3.10 14.50 3.78 15.58 3.78 15.58 4.10
                 12.78 4.10 12.78 1.96 10.30 1.96 10.30 3.78 11.38 3.78
                 11.38 3.16 11.70 3.16 11.70 3.78 12.78 3.78 12.78 4.10
                 9.98 4.10 9.98 1.96 7.50 1.96 7.50 3.78 8.58 3.78 8.58 3.10
                 8.90 3.10 8.90 3.78 9.98 3.78 9.98 4.10 7.18 4.10 7.18 1.96
                 4.70 1.96 4.70 3.78 5.78 3.78 5.78 3.16 6.10 3.16 6.10 3.78
                 7.18 3.78 7.18 4.10 4.38 4.10 4.38 1.96 1.90 1.96 1.90 3.78
                 2.98 3.78 2.98 3.10 3.30 3.10 3.30 3.78 4.38 3.78 4.38 4.10
                 0.18 4.10 0.18 3.16 0.50 3.16 0.50 3.78 1.58 3.78 1.58 1.96
                 0.18 1.96 0.18 1.64 22.90 1.64 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  23.68 0.90 22.20 0.90 22.20 1.32 21.88 1.32 21.88 0.90
                 20.80 0.90 20.80 1.32 20.48 1.32 20.48 0.90 19.40 0.90
                 19.40 1.32 19.08 1.32 19.08 0.90 18.00 0.90 18.00 1.32
                 17.68 1.32 17.68 0.90 16.60 0.90 16.60 1.32 16.28 1.32
                 16.28 0.90 15.20 0.90 15.20 1.32 14.88 1.32 14.88 0.90
                 13.80 0.90 13.80 1.32 13.48 1.32 13.48 0.90 12.40 0.90
                 12.40 1.32 12.08 1.32 12.08 0.90 11.00 0.90 11.00 1.32
                 10.68 1.32 10.68 0.90 9.60 0.90 9.60 1.32 9.28 1.32 9.28 0.90
                 8.20 0.90 8.20 1.32 7.88 1.32 7.88 0.90 6.80 0.90 6.80 1.32
                 6.48 1.32 6.48 0.90 5.40 0.90 5.40 1.32 5.08 1.32 5.08 0.90
                 4.00 0.90 4.00 1.32 3.68 1.32 3.68 0.90 2.60 0.90 2.60 1.32
                 2.28 1.32 2.28 0.90 1.20 0.90 1.20 1.32 0.88 1.32 0.88 0.90
                 0.00 0.90 0.00 -0.90 23.68 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  23.68 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.42 1.20 4.42
                 1.20 4.86 2.28 4.86 2.28 4.42 2.60 4.42 2.60 4.86 3.68 4.86
                 3.68 4.42 4.00 4.42 4.00 4.86 5.08 4.86 5.08 4.42 5.40 4.42
                 5.40 4.86 6.48 4.86 6.48 4.42 6.80 4.42 6.80 4.86 7.88 4.86
                 7.88 4.42 8.20 4.42 8.20 4.86 9.28 4.86 9.28 4.42 9.60 4.42
                 9.60 4.86 10.68 4.86 10.68 4.42 11.00 4.42 11.00 4.86
                 12.08 4.86 12.08 4.42 12.40 4.42 12.40 4.86 13.48 4.86
                 13.48 4.42 13.80 4.42 13.80 4.86 14.88 4.86 14.88 4.42
                 15.20 4.42 15.20 4.86 16.28 4.86 16.28 4.42 16.60 4.42
                 16.60 4.86 17.68 4.86 17.68 4.42 18.00 4.42 18.00 4.86
                 19.08 4.86 19.08 4.42 19.40 4.42 19.40 4.86 20.48 4.86
                 20.48 4.42 20.80 4.42 20.80 4.86 21.88 4.86 21.88 4.42
                 22.20 4.42 22.20 4.86 23.68 4.86 ;
        END
    END vdd!
END inv_64

MACRO inv_6
    CLASS CORE ;
    FOREIGN inv_6 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.20 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.04  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.34 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.90 4.20 1.58 4.20 1.58 3.70 0.50 3.70 0.50 4.20 0.18 4.20
                 0.18 3.16 0.50 3.16 0.50 3.38 1.58 3.38 1.58 3.04 1.44 3.04
                 1.44 2.72 1.58 2.72 1.58 1.96 0.18 1.96 0.18 1.64 1.90 1.64 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  3.20 0.90 2.60 0.90 2.60 2.18 2.28 2.18 2.28 0.90 1.20 0.90
                 1.20 1.32 0.88 1.32 0.88 0.90 0.00 0.90 0.00 -0.90 3.20 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  3.20 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.34 1.20 4.34
                 1.20 4.86 2.28 4.86 2.28 3.10 2.60 3.10 2.60 4.86 3.20 4.86 ;
        END
    END vdd!
END inv_6

MACRO inv_48
    CLASS CORE ;
    FOREIGN inv_48 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 17.92 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 16.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.34 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 24.95  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  17.30 1.96 15.90 1.96 15.90 3.38 16.98 3.38 16.98 3.16
                 17.30 3.16 17.30 4.20 16.98 4.20 16.98 3.70 15.90 3.70
                 15.90 4.20 15.58 4.20 15.58 3.04 15.52 3.04 15.52 2.72
                 15.58 2.72 15.58 1.96 14.50 1.96 14.50 3.38 15.58 3.38
                 15.58 3.70 14.50 3.70 14.50 4.20 14.18 4.20 14.18 1.96
                 11.70 1.96 11.70 3.38 12.78 3.38 12.78 3.16 13.10 3.16
                 13.10 3.38 14.18 3.38 14.18 3.70 13.10 3.70 13.10 4.20
                 12.78 4.20 12.78 3.70 11.70 3.70 11.70 4.20 11.38 4.20
                 11.38 1.96 10.30 1.96 10.30 3.38 11.38 3.38 11.38 3.70
                 10.30 3.70 10.30 4.20 9.98 4.20 9.98 1.96 7.50 1.96 7.50 3.38
                 8.58 3.38 8.58 3.16 8.90 3.16 8.90 3.38 9.98 3.38 9.98 3.70
                 8.90 3.70 8.90 4.20 8.58 4.20 8.58 3.70 7.50 3.70 7.50 4.20
                 7.18 4.20 7.18 1.96 6.10 1.96 6.10 3.38 7.18 3.38 7.18 3.70
                 6.10 3.70 6.10 4.20 5.78 4.20 5.78 1.96 3.30 1.96 3.30 3.38
                 4.38 3.38 4.38 3.16 4.70 3.16 4.70 3.38 5.78 3.38 5.78 3.70
                 4.70 3.70 4.70 4.20 4.38 4.20 4.38 3.70 3.30 3.70 3.30 4.20
                 2.98 4.20 2.98 1.96 1.90 1.96 1.90 3.38 2.98 3.38 2.98 3.70
                 1.90 3.70 1.90 4.20 1.58 4.20 1.58 3.70 0.50 3.70 0.50 4.20
                 0.18 4.20 0.18 3.16 0.50 3.16 0.50 3.38 1.58 3.38 1.58 1.96
                 0.18 1.96 0.18 1.64 17.30 1.64 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  17.92 0.90 16.60 0.90 16.60 1.32 16.28 1.32 16.28 0.90
                 15.20 0.90 15.20 1.32 14.88 1.32 14.88 0.90 13.80 0.90
                 13.80 1.32 13.48 1.32 13.48 0.90 12.40 0.90 12.40 1.32
                 12.08 1.32 12.08 0.90 11.00 0.90 11.00 1.32 10.68 1.32
                 10.68 0.90 9.60 0.90 9.60 1.32 9.28 1.32 9.28 0.90 8.20 0.90
                 8.20 1.32 7.88 1.32 7.88 0.90 6.80 0.90 6.80 1.32 6.48 1.32
                 6.48 0.90 5.40 0.90 5.40 1.32 5.08 1.32 5.08 0.90 4.00 0.90
                 4.00 1.32 3.68 1.32 3.68 0.90 2.60 0.90 2.60 1.32 2.28 1.32
                 2.28 0.90 1.20 0.90 1.20 1.32 0.88 1.32 0.88 0.90 0.00 0.90
                 0.00 -0.90 17.92 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  17.92 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.34 1.20 4.34
                 1.20 4.86 2.28 4.86 2.28 4.34 2.60 4.34 2.60 4.86 3.68 4.86
                 3.68 4.34 4.00 4.34 4.00 4.86 5.08 4.86 5.08 4.34 5.40 4.34
                 5.40 4.86 6.48 4.86 6.48 4.34 6.80 4.34 6.80 4.86 7.88 4.86
                 7.88 4.34 8.20 4.34 8.20 4.86 9.28 4.86 9.28 4.34 9.60 4.34
                 9.60 4.86 10.68 4.86 10.68 4.34 11.00 4.34 11.00 4.86
                 12.08 4.86 12.08 4.34 12.40 4.34 12.40 4.86 13.48 4.86
                 13.48 4.34 13.80 4.34 13.80 4.86 14.88 4.86 14.88 4.34
                 15.20 4.34 15.20 4.86 16.28 4.86 16.28 4.34 16.60 4.34
                 16.60 4.86 17.92 4.86 ;
        END
    END vdd!
END inv_48

MACRO inv_4
    CLASS CORE ;
    FOREIGN inv_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.56 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.34 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.90 4.14 1.58 4.14 1.58 3.86 0.50 3.86 0.50 4.14 0.18 4.14
                 0.18 3.26 0.50 3.26 0.50 3.54 1.58 3.54 1.58 3.04 1.44 3.04
                 1.44 2.72 1.58 2.72 1.58 1.96 0.18 1.96 0.18 1.64 1.90 1.64 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  2.56 0.90 1.20 0.90 1.20 1.32 0.88 1.32 0.88 0.90 0.00 0.90
                 0.00 -0.90 2.56 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  2.56 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.42 1.20 4.42
                 1.20 4.86 2.56 4.86 ;
        END
    END vdd!
END inv_4

MACRO inv_32
    CLASS CORE ;
    FOREIGN inv_32 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.16 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 10.89  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.34 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 17.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  11.70 1.96 10.30 1.96 10.30 3.78 11.38 3.78 11.38 3.16
                 11.70 3.16 11.70 4.10 9.98 4.10 9.98 3.04 9.76 3.04 9.76 2.72
                 9.98 2.72 9.98 1.96 7.50 1.96 7.50 3.78 8.58 3.78 8.58 3.10
                 8.90 3.10 8.90 3.78 9.98 3.78 9.98 4.10 7.18 4.10 7.18 1.96
                 4.70 1.96 4.70 3.78 5.78 3.78 5.78 3.16 6.10 3.16 6.10 3.78
                 7.18 3.78 7.18 4.10 4.38 4.10 4.38 1.96 1.90 1.96 1.90 3.78
                 2.98 3.78 2.98 3.10 3.30 3.10 3.30 3.78 4.38 3.78 4.38 4.10
                 0.18 4.10 0.18 3.16 0.50 3.16 0.50 3.78 1.58 3.78 1.58 1.96
                 0.18 1.96 0.18 1.64 11.70 1.64 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  12.16 0.90 11.00 0.90 11.00 1.32 10.68 1.32 10.68 0.90
                 9.60 0.90 9.60 1.32 9.28 1.32 9.28 0.90 8.20 0.90 8.20 1.32
                 7.88 1.32 7.88 0.90 6.80 0.90 6.80 1.32 6.48 1.32 6.48 0.90
                 5.40 0.90 5.40 1.32 5.08 1.32 5.08 0.90 4.00 0.90 4.00 1.32
                 3.68 1.32 3.68 0.90 2.60 0.90 2.60 1.32 2.28 1.32 2.28 0.90
                 1.20 0.90 1.20 1.32 0.88 1.32 0.88 0.90 0.00 0.90 0.00 -0.90
                 12.16 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  12.16 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.42 1.20 4.42
                 1.20 4.86 2.28 4.86 2.28 4.42 2.60 4.42 2.60 4.86 3.68 4.86
                 3.68 4.42 4.00 4.42 4.00 4.86 5.08 4.86 5.08 4.42 5.40 4.42
                 5.40 4.86 6.48 4.86 6.48 4.42 6.80 4.42 6.80 4.86 7.88 4.86
                 7.88 4.42 8.20 4.42 8.20 4.86 9.28 4.86 9.28 4.42 9.60 4.42
                 9.60 4.86 10.68 4.86 10.68 4.42 11.00 4.42 11.00 4.86
                 12.16 4.86 ;
        END
    END vdd!
END inv_32

MACRO inv_3
    CLASS CORE ;
    FOREIGN inv_3 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.20 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.47  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.34 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.61  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.90 4.34 0.18 4.34 0.18 4.02 1.58 4.02 1.58 3.04 1.44 3.04
                 1.44 2.72 1.58 2.72 1.58 1.66 0.18 1.66 0.18 1.34 1.90 1.34 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  3.20 0.90 2.60 0.90 2.60 1.76 2.28 1.76 2.28 0.90 1.20 0.90
                 1.20 1.00 0.88 1.00 0.88 0.90 0.00 0.90 0.00 -0.90 3.20 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  3.20 6.66 0.00 6.66 0.00 4.86 2.28 4.86 2.28 4.30 2.60 4.30
                 2.60 4.86 3.20 4.86 ;
        END
    END vdd!
END inv_3

MACRO inv_24
    CLASS CORE ;
    FOREIGN inv_24 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.60 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 8.16  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.34 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 13.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.90 1.96 7.50 1.96 7.50 2.72 7.52 2.72 7.52 3.04 7.50 3.04
                 7.50 3.38 8.58 3.38 8.58 3.16 8.90 3.16 8.90 4.20 8.58 4.20
                 8.58 3.70 7.50 3.70 7.50 4.20 7.18 4.20 7.18 1.96 6.10 1.96
                 6.10 3.38 7.18 3.38 7.18 3.70 6.10 3.70 6.10 4.20 5.78 4.20
                 5.78 1.96 3.30 1.96 3.30 3.38 4.38 3.38 4.38 3.16 4.70 3.16
                 4.70 3.38 5.78 3.38 5.78 3.70 4.70 3.70 4.70 4.20 4.38 4.20
                 4.38 3.70 3.30 3.70 3.30 4.20 2.98 4.20 2.98 1.96 1.90 1.96
                 1.90 3.38 2.98 3.38 2.98 3.70 1.90 3.70 1.90 4.20 1.58 4.20
                 1.58 3.70 0.50 3.70 0.50 4.20 0.18 4.20 0.18 3.16 0.50 3.16
                 0.50 3.38 1.58 3.38 1.58 1.96 0.18 1.96 0.18 1.64 8.90 1.64 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  9.60 0.90 8.20 0.90 8.20 1.32 7.88 1.32 7.88 0.90 6.80 0.90
                 6.80 1.32 6.48 1.32 6.48 0.90 5.40 0.90 5.40 1.32 5.08 1.32
                 5.08 0.90 4.00 0.90 4.00 1.32 3.68 1.32 3.68 0.90 2.60 0.90
                 2.60 1.32 2.28 1.32 2.28 0.90 1.20 0.90 1.20 1.32 0.88 1.32
                 0.88 0.90 0.00 0.90 0.00 -0.90 9.60 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  9.60 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.34 1.20 4.34
                 1.20 4.86 2.28 4.86 2.28 4.34 2.60 4.34 2.60 4.86 3.68 4.86
                 3.68 4.34 4.00 4.34 4.00 4.86 5.08 4.86 5.08 4.34 5.40 4.34
                 5.40 4.86 6.48 4.86 6.48 4.34 6.80 4.34 6.80 4.86 7.88 4.86
                 7.88 4.34 8.20 4.34 8.20 4.86 9.60 4.86 ;
        END
    END vdd!
END inv_24

MACRO inv_20
    CLASS CORE ;
    FOREIGN inv_20 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 6.80  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.34 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 11.19  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.50 1.96 6.10 1.96 6.10 2.72 6.24 2.72 6.24 3.04 6.10 3.04
                 6.10 3.58 7.50 3.58 7.50 4.54 7.18 4.54 7.18 3.90 6.10 3.90
                 6.10 4.54 5.78 4.54 5.78 1.96 1.90 1.96 1.90 3.58 5.78 3.58
                 5.78 3.90 4.70 3.90 4.70 4.54 4.38 4.54 4.38 3.90 3.30 3.90
                 3.30 4.54 2.98 4.54 2.98 3.90 1.90 3.90 1.90 4.54 1.58 4.54
                 1.58 3.90 0.50 3.90 0.50 4.54 0.18 4.54 0.18 3.58 1.58 3.58
                 1.58 1.96 0.18 1.96 0.18 1.64 7.50 1.64 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 0.90 6.80 0.90 6.80 1.32 6.48 1.32 6.48 0.90 5.40 0.90
                 5.40 1.32 5.08 1.32 5.08 0.90 4.00 0.90 4.00 1.32 3.68 1.32
                 3.68 0.90 2.60 0.90 2.60 1.32 2.28 1.32 2.28 0.90 1.20 0.90
                 1.20 1.32 0.88 1.32 0.88 0.90 0.00 0.90 0.00 -0.90 7.68 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 2.28 4.86 2.28 4.22 2.60 4.22 2.60 4.86 3.68 4.86
                 3.68 4.22 4.00 4.22 4.00 4.86 5.08 4.86 5.08 4.22 5.40 4.22
                 5.40 4.86 6.48 4.86 6.48 4.22 6.80 4.22 6.80 4.86 7.68 4.86 ;
        END
    END vdd!
END inv_20

MACRO inv_2
    CLASS CORE ;
    FOREIGN inv_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 1.92 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.48 2.08 1.12 2.66 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.76 3.58 1.44 3.58 1.44 4.54 1.12 4.54 1.12 3.26 1.44 3.26
                 1.44 1.70 1.12 1.70 1.12 1.38 1.76 1.38 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  1.92 0.90 0.74 0.90 0.74 1.32 0.42 1.32 0.42 0.90 0.00 0.90
                 0.00 -0.90 1.92 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  1.92 6.66 0.00 6.66 0.00 4.86 0.42 4.86 0.42 3.56 0.74 3.56
                 0.74 4.86 1.92 4.86 ;
        END
    END vdd!
END inv_2

MACRO inv_16
    CLASS CORE ;
    FOREIGN inv_16 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 5.44  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.34 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 9.22  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  6.10 1.96 4.70 1.96 4.70 2.72 4.96 2.72 4.96 3.04 4.70 3.04
                 4.70 3.78 5.78 3.78 5.78 3.16 6.10 3.16 6.10 4.10 4.38 4.10
                 4.38 1.96 1.90 1.96 1.90 3.78 2.98 3.78 2.98 3.10 3.30 3.10
                 3.30 3.78 4.38 3.78 4.38 4.10 0.18 4.10 0.18 3.16 0.50 3.16
                 0.50 3.78 1.58 3.78 1.58 1.96 0.18 1.96 0.18 1.64 6.10 1.64 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 0.90 5.40 0.90 5.40 1.32 5.08 1.32 5.08 0.90 4.00 0.90
                 4.00 1.32 3.68 1.32 3.68 0.90 2.60 0.90 2.60 1.32 2.28 1.32
                 2.28 0.90 1.20 0.90 1.20 1.32 0.88 1.32 0.88 0.90 0.00 0.90
                 0.00 -0.90 6.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.42 1.20 4.42
                 1.20 4.86 2.28 4.86 2.28 4.42 2.60 4.42 2.60 4.86 3.68 4.86
                 3.68 4.42 4.00 4.42 4.00 4.86 5.08 4.86 5.08 4.42 5.40 4.42
                 5.40 4.86 6.40 4.86 ;
        END
    END vdd!
END inv_16

MACRO inv_12
    CLASS CORE ;
    FOREIGN inv_12 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 7.26  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.70 1.96 3.30 1.96 3.30 2.72 3.68 2.72 3.68 3.04 3.30 3.04
                 3.30 3.38 4.38 3.38 4.38 3.16 4.70 3.16 4.70 4.20 4.38 4.20
                 4.38 3.70 3.30 3.70 3.30 4.20 2.98 4.20 2.98 1.96 1.90 1.96
                 1.90 3.38 2.98 3.38 2.98 3.70 1.90 3.70 1.90 4.20 1.58 4.20
                 1.58 3.70 0.50 3.70 0.50 4.20 0.18 4.20 0.18 3.16 0.50 3.16
                 0.50 3.38 1.58 3.38 1.58 1.96 0.18 1.96 0.18 1.64 4.70 1.64 ;
        END
    END x
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 4.08  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.34 1.12 3.04 ;
        END
    END a
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.34 1.20 4.34
                 1.20 4.86 2.28 4.86 2.28 4.34 2.60 4.34 2.60 4.86 3.68 4.86
                 3.68 4.34 4.00 4.34 4.00 4.86 5.12 4.86 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 0.90 4.00 0.90 4.00 1.32 3.68 1.32 3.68 0.90 2.60 0.90
                 2.60 1.32 2.28 1.32 2.28 0.90 1.20 0.90 1.20 1.32 0.88 1.32
                 0.88 0.90 0.00 0.90 0.00 -0.90 5.12 -0.90 ;
        END
    END gnd!
END inv_12

MACRO inv_10
    CLASS CORE ;
    FOREIGN inv_10 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.48 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.40  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.34 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.59  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.30 1.96 1.90 1.96 1.90 3.58 3.30 3.58 3.30 4.54 2.98 4.54
                 2.98 3.90 1.90 3.90 1.90 4.54 1.58 4.54 1.58 3.90 0.50 3.90
                 0.50 4.54 0.18 4.54 0.18 3.58 1.58 3.58 1.58 3.04 1.44 3.04
                 1.44 2.72 1.58 2.72 1.58 1.96 0.18 1.96 0.18 1.64 3.30 1.64 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  4.48 0.90 4.00 0.90 4.00 2.18 3.68 2.18 3.68 0.90 2.60 0.90
                 2.60 1.32 2.28 1.32 2.28 0.90 1.20 0.90 1.20 1.32 0.88 1.32
                 0.88 0.90 0.00 0.90 0.00 -0.90 4.48 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  4.48 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 2.28 4.86 2.28 4.22 2.60 4.22 2.60 4.86 3.68 4.86
                 3.68 3.10 4.00 3.10 4.00 4.86 4.48 4.86 ;
        END
    END vdd!
END inv_10

MACRO inv_1
    CLASS CORE ;
    FOREIGN inv_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 1.92 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.48 2.62 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.76 3.78 1.44 3.78 1.44 4.34 1.12 4.34 1.12 3.46 1.44 3.46
                 1.44 1.70 1.12 1.70 1.12 1.38 1.76 1.38 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  1.92 0.90 0.74 0.90 0.74 1.32 0.42 1.32 0.42 0.90 0.00 0.90
                 0.00 -0.90 1.92 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  1.92 6.66 0.00 6.66 0.00 4.86 0.42 4.86 0.42 3.56 0.74 3.56
                 0.74 4.86 1.92 4.86 ;
        END
    END vdd!
END inv_1

MACRO inv_0
    CLASS CORE ;
    FOREIGN inv_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 1.92 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.45  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.48 2.62 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.76 3.78 1.44 3.78 1.44 4.34 1.12 4.34 1.12 3.46 1.44 3.46
                 1.44 1.70 1.12 1.70 1.12 1.38 1.76 1.38 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  1.92 0.90 0.74 0.90 0.74 1.32 0.42 1.32 0.42 0.90 0.00 0.90
                 0.00 -0.90 1.92 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  1.92 6.66 0.00 6.66 0.00 4.86 0.42 4.86 0.42 3.56 0.74 3.56
                 0.74 4.86 1.92 4.86 ;
        END
    END vdd!
END inv_0

MACRO gclklatp_8
    CLASS CORE ;
    FOREIGN gclklatp_8 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.75  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.40 2.08 10.72 2.82 ;
        END
    END ck
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END g
    PIN gck
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 8.05  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  21.72 4.46 21.40 4.46 21.40 3.80 20.32 3.80 20.32 4.46
                 20.00 4.46 20.00 3.80 18.92 3.80 18.92 4.46 18.60 4.46
                 18.60 3.80 17.52 3.80 17.52 4.46 17.20 4.46 17.20 3.80
                 16.12 3.80 16.12 4.46 15.80 4.46 15.80 3.48 21.40 3.48
                 21.40 3.04 21.28 3.04 21.28 2.72 21.40 2.72 21.40 1.62
                 15.80 1.62 15.80 1.30 21.72 1.30 ;
        END
    END gck
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  22.40 0.90 1.20 0.90 1.20 1.30 0.88 1.30 0.88 0.90 0.00 0.90
                 0.00 -0.90 22.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  22.40 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.16 1.20 4.16
                 1.20 4.86 4.53 4.86 4.53 4.62 4.85 4.62 4.85 4.86 9.83 4.86
                 9.83 4.00 10.15 4.00 10.15 4.86 11.23 4.86 11.23 4.00
                 11.55 4.00 11.55 4.86 12.66 4.86 12.66 4.00 12.98 4.00
                 12.98 4.86 14.06 4.86 14.06 4.00 14.38 4.00 14.38 4.86
                 16.50 4.86 16.50 4.37 16.82 4.37 16.82 4.86 17.90 4.86
                 17.90 4.37 18.22 4.37 18.22 4.86 19.30 4.86 19.30 4.37
                 19.62 4.37 19.62 4.86 20.70 4.86 20.70 4.37 21.02 4.37
                 21.02 4.86 22.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  17.20 2.68 14.73 2.68 14.73 3.36 15.08 3.36 15.08 4.54
                 14.76 4.54 14.76 3.68 13.68 3.68 13.68 4.54 13.36 4.54
                 13.36 3.68 12.25 3.68 12.25 4.54 11.93 4.54 11.93 3.68
                 10.85 3.68 10.85 4.54 10.53 4.54 10.53 3.68 9.45 3.68
                 9.45 4.54 9.13 4.54 9.13 3.68 9.12 3.68 9.12 3.36 14.41 3.36
                 14.41 2.18 13.01 2.18 13.01 1.86 14.73 1.86 14.73 2.36
                 17.20 2.36 ;
        RECT  8.82 1.22 15.43 1.54 ;
        POLYGON  8.77 4.03 8.45 4.03 8.45 2.50 7.06 2.50 7.06 2.62 5.28 2.62
                 5.28 2.30 6.74 2.30 6.74 2.18 8.15 2.18 8.15 1.88 8.47 1.88
                 8.47 2.18 8.77 2.18 ;
        POLYGON  7.84 4.54 5.17 4.54 5.17 3.90 2.58 3.90 2.58 4.54 2.26 4.54
                 2.26 1.28 2.58 1.28 2.58 3.58 5.49 3.58 5.49 4.22 7.52 4.22
                 7.52 2.82 7.84 2.82 ;
        POLYGON  7.12 3.90 5.82 3.90 5.82 3.58 6.80 3.58 6.80 2.94 7.12 2.94 ;
        RECT  6.02 1.52 6.90 1.86 ;
        POLYGON  5.78 3.26 4.38 3.26 4.38 2.62 3.58 2.62 3.58 2.30 4.38 2.30
                 4.38 1.65 5.70 1.65 5.70 1.97 4.70 1.97 4.70 2.94 5.78 2.94 ;
        RECT  3.05 1.26 4.06 1.58 ;
        RECT  2.96 4.22 4.06 4.54 ;
        POLYGON  1.88 1.94 0.18 1.94 0.18 1.44 0.50 1.44 0.50 1.62 1.56 1.62
                 1.56 1.38 1.88 1.38 ;
        POLYGON  1.88 4.54 1.56 4.54 1.56 3.76 0.50 3.76 0.50 4.48 0.18 4.48
                 0.18 3.44 1.88 3.44 ;
    END
END gclklatp_8

MACRO gclklatp_4
    CLASS CORE ;
    FOREIGN gclklatp_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.64 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.62  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  9.76 2.08 10.08 2.82 ;
        END
    END ck
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END g
    PIN gck
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.62  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.11 4.46 15.79 4.46 15.79 3.80 14.71 3.80 14.71 4.46
                 14.39 4.46 14.39 3.80 13.31 3.80 13.31 4.46 12.99 4.46
                 12.99 3.48 15.79 3.48 15.79 3.04 15.52 3.04 15.52 2.72
                 15.79 2.72 15.79 1.62 12.99 1.62 12.99 1.30 16.11 1.30 ;
        END
    END gck
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 0.90 1.20 0.90 1.20 1.30 0.88 1.30 0.88 0.90 0.00 0.90
                 0.00 -0.90 16.64 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.16 1.20 4.16
                 1.20 4.86 4.53 4.86 4.53 4.62 4.85 4.62 4.85 4.86 9.83 4.86
                 9.83 4.00 10.15 4.00 10.15 4.86 11.26 4.86 11.26 4.00
                 11.58 4.00 11.58 4.86 13.69 4.86 13.69 4.37 14.01 4.37
                 14.01 4.86 15.09 4.86 15.09 4.37 15.41 4.37 15.41 4.86
                 16.64 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  14.53 2.68 12.27 2.68 12.27 3.36 12.28 3.36 12.28 4.54
                 11.96 4.54 11.96 3.68 10.85 3.68 10.85 4.54 10.53 4.54
                 10.53 3.68 9.45 3.68 9.45 4.54 9.13 4.54 9.13 3.36 11.95 3.36
                 11.95 2.18 11.61 2.18 11.61 1.86 12.27 1.86 12.27 2.36
                 14.53 2.36 ;
        RECT  8.83 1.22 12.63 1.54 ;
        POLYGON  8.77 4.03 8.45 4.03 8.45 2.50 7.06 2.50 7.06 2.62 5.28 2.62
                 5.28 2.30 6.74 2.30 6.74 2.18 8.15 2.18 8.15 1.88 8.47 1.88
                 8.47 2.18 8.77 2.18 ;
        POLYGON  7.84 4.54 5.17 4.54 5.17 3.90 2.58 3.90 2.58 4.54 2.26 4.54
                 2.26 1.28 2.58 1.28 2.58 3.58 5.49 3.58 5.49 4.22 7.52 4.22
                 7.52 2.82 7.84 2.82 ;
        POLYGON  7.12 3.90 5.82 3.90 5.82 3.58 6.80 3.58 6.80 2.94 7.12 2.94 ;
        RECT  6.02 1.52 6.90 1.86 ;
        POLYGON  5.78 3.26 4.38 3.26 4.38 2.62 3.58 2.62 3.58 2.30 4.38 2.30
                 4.38 1.65 5.70 1.65 5.70 1.97 4.70 1.97 4.70 2.94 5.78 2.94 ;
        RECT  3.05 1.26 4.06 1.58 ;
        RECT  2.96 4.22 4.06 4.54 ;
        POLYGON  1.88 1.94 0.18 1.94 0.18 1.44 0.50 1.44 0.50 1.62 1.56 1.62
                 1.56 1.38 1.88 1.38 ;
        POLYGON  1.88 4.54 1.56 4.54 1.56 3.76 0.50 3.76 0.50 4.48 0.18 4.48
                 0.18 3.44 1.88 3.44 ;
    END
END gclklatp_4

MACRO gclklatp_2
    CLASS CORE ;
    FOREIGN gclklatp_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.36 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.62  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  9.76 2.08 10.08 2.82 ;
        END
    END ck
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END g
    PIN gck
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.92  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  15.20 3.80 14.71 3.80 14.71 4.46 14.39 4.46 14.39 3.80
                 13.31 3.80 13.31 4.46 12.99 4.46 12.99 3.48 14.88 3.48
                 14.88 1.64 12.99 1.64 12.99 1.32 15.20 1.32 ;
        END
    END gck
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  15.36 0.90 1.20 0.90 1.20 1.30 0.88 1.30 0.88 0.90 0.00 0.90
                 0.00 -0.90 15.36 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  15.36 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.16 1.20 4.16
                 1.20 4.86 4.53 4.86 4.53 4.62 4.85 4.62 4.85 4.86 9.83 4.86
                 9.83 4.00 10.15 4.00 10.15 4.86 11.26 4.86 11.26 4.00
                 11.58 4.00 11.58 4.86 13.69 4.86 13.69 4.37 14.01 4.37
                 14.01 4.86 15.36 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  13.74 2.68 12.27 2.68 12.27 3.36 12.28 3.36 12.28 4.54
                 11.96 4.54 11.96 3.68 10.85 3.68 10.85 4.54 10.53 4.54
                 10.53 3.68 9.45 3.68 9.45 4.54 9.13 4.54 9.13 3.36 11.95 3.36
                 11.95 2.18 11.61 2.18 11.61 1.86 12.27 1.86 12.27 2.36
                 13.74 2.36 ;
        RECT  8.83 1.22 12.63 1.54 ;
        POLYGON  8.77 4.03 8.45 4.03 8.45 2.50 7.06 2.50 7.06 2.62 5.28 2.62
                 5.28 2.30 6.74 2.30 6.74 2.18 8.15 2.18 8.15 1.88 8.47 1.88
                 8.47 2.18 8.77 2.18 ;
        POLYGON  7.84 4.54 5.17 4.54 5.17 3.90 2.58 3.90 2.58 4.54 2.26 4.54
                 2.26 1.28 2.58 1.28 2.58 3.58 5.49 3.58 5.49 4.22 7.52 4.22
                 7.52 2.82 7.84 2.82 ;
        POLYGON  7.12 3.90 5.82 3.90 5.82 3.58 6.80 3.58 6.80 2.94 7.12 2.94 ;
        RECT  6.02 1.52 6.90 1.86 ;
        POLYGON  5.78 3.26 4.38 3.26 4.38 2.62 3.58 2.62 3.58 2.30 4.38 2.30
                 4.38 1.65 5.70 1.65 5.70 1.97 4.70 1.97 4.70 2.94 5.78 2.94 ;
        RECT  3.05 1.26 4.06 1.58 ;
        RECT  2.96 4.22 4.06 4.54 ;
        POLYGON  1.88 1.94 0.18 1.94 0.18 1.44 0.50 1.44 0.50 1.62 1.56 1.62
                 1.56 1.38 1.88 1.38 ;
        POLYGON  1.88 4.54 1.56 4.54 1.56 3.76 0.50 3.76 0.50 4.48 0.18 4.48
                 0.18 3.44 1.88 3.44 ;
    END
END gclklatp_2

MACRO gclklatp_1
    CLASS CORE ;
    FOREIGN gclklatp_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.80 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.44 3.04 8.57 3.04 8.57 1.65 8.46 1.54 6.00 1.54 6.00 1.22
                 8.60 1.22 8.89 1.51 8.89 2.72 9.44 2.72 ;
        END
    END ck
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END g
    PIN gck
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.46  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.64 3.04 12.46 3.04 12.46 3.80 11.64 3.80 11.64 4.44
                 11.32 4.44 11.32 3.48 12.14 3.48 12.14 1.64 12.10 1.64
                 12.10 1.32 12.46 1.32 12.46 2.72 12.64 2.72 ;
        END
    END gck
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  12.80 0.90 11.72 0.90 11.72 1.32 11.40 1.32 11.40 0.90
                 1.20 0.90 1.20 1.30 0.88 1.30 0.88 0.90 0.00 0.90 0.00 -0.90
                 12.80 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  12.80 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.16 1.20 4.16
                 1.20 4.86 4.53 4.86 4.53 4.62 4.85 4.62 4.85 4.86 8.61 4.86
                 8.61 4.00 8.93 4.00 8.93 4.86 10.04 4.86 10.04 4.00 10.36 4.00
                 10.36 4.86 12.02 4.86 12.02 4.12 12.34 4.12 12.34 4.86
                 12.80 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  11.01 3.03 10.56 3.03 10.56 3.68 9.63 3.68 9.63 4.54 9.31 4.54
                 9.31 3.36 10.22 3.36 10.22 2.71 10.69 2.71 10.69 1.64
                 11.01 1.64 ;
        POLYGON  10.31 1.54 9.63 1.54 9.63 1.96 9.31 1.96 9.31 1.22 10.31 1.22 ;
        POLYGON  8.25 4.54 5.82 4.54 5.82 4.22 7.93 4.22 7.93 1.88 8.25 1.88 ;
        POLYGON  7.54 2.92 7.46 2.92 7.46 3.90 2.58 3.90 2.58 4.54 2.26 4.54
                 2.26 1.28 2.58 1.28 2.58 3.58 7.14 3.58 7.14 2.60 7.54 2.60 ;
        POLYGON  6.68 3.26 6.28 3.26 6.28 2.94 6.36 2.94 6.36 2.62 5.26 2.62
                 5.26 2.30 6.36 2.30 6.36 1.88 6.68 1.88 ;
        POLYGON  5.78 3.26 4.38 3.26 4.38 2.62 3.58 2.62 3.58 2.30 4.38 2.30
                 4.38 1.66 5.70 1.66 5.70 1.98 4.70 1.98 4.70 2.94 5.78 2.94 ;
        RECT  3.05 1.26 4.06 1.58 ;
        RECT  2.96 4.22 4.06 4.54 ;
        POLYGON  1.88 1.94 0.18 1.94 0.18 1.44 0.50 1.44 0.50 1.62 1.56 1.62
                 1.56 1.38 1.88 1.38 ;
        POLYGON  1.88 4.54 1.56 4.54 1.56 3.76 0.50 3.76 0.50 4.48 0.18 4.48
                 0.18 3.44 1.88 3.44 ;
    END
END gclklatp_1

MACRO gclklatn_8
    CLASS CORE ;
    FOREIGN gclklatn_8 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.76 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  11.48 2.40 11.04 2.40 11.04 2.26 8.59 2.26 8.59 1.54 6.02 1.54
                 6.02 1.22 8.91 1.22 8.91 1.94 11.48 1.94 ;
        END
    END ck
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END g
    PIN gck
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 8.34  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  21.54 4.44 21.22 4.44 21.22 1.63 18.74 1.63 18.74 3.36
                 21.22 3.36 21.22 3.68 20.14 3.68 20.14 4.44 19.82 4.44
                 19.82 3.68 18.74 3.68 18.74 4.44 18.42 4.44 18.42 3.68
                 17.34 3.68 17.34 4.44 17.02 4.44 17.02 3.68 15.94 3.68
                 15.94 4.44 15.62 4.44 15.62 3.36 18.42 3.36 18.42 1.63
                 15.61 1.63 15.61 1.31 21.54 1.31 ;
        END
    END gck
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.76 0.90 1.20 0.90 1.20 1.30 0.88 1.30 0.88 0.90 0.00 0.90
                 0.00 -0.90 21.76 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.76 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.13 1.20 4.13
                 1.20 4.86 4.53 4.86 4.53 4.60 4.85 4.60 4.85 4.86 9.33 4.86
                 9.33 3.99 9.65 3.99 9.65 4.86 10.73 4.86 10.73 3.99 11.05 3.99
                 11.05 4.86 16.32 4.86 16.32 4.11 16.64 4.11 16.64 4.86
                 17.72 4.86 17.72 4.12 18.04 4.12 18.04 4.86 19.12 4.86
                 19.12 4.11 19.44 4.11 19.44 4.86 20.52 4.86 20.52 4.11
                 20.84 4.11 20.84 4.86 21.76 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  17.37 2.58 15.26 2.58 15.26 4.54 14.94 4.54 14.94 3.30
                 13.86 3.30 13.86 3.90 13.54 3.90 13.54 3.30 12.43 3.30
                 12.43 3.88 12.11 3.88 12.11 2.82 12.43 2.82 12.43 2.98
                 14.94 2.98 14.94 1.54 9.25 1.54 9.25 1.22 15.26 1.22
                 15.26 2.26 17.37 2.26 ;
        POLYGON  14.56 4.54 11.43 4.54 11.43 3.30 10.35 3.30 10.35 4.54
                 10.03 4.54 10.03 3.30 8.95 3.30 8.95 4.54 8.63 4.54 8.63 2.98
                 11.75 2.98 11.75 4.22 12.84 4.22 12.84 3.62 13.16 3.62
                 13.16 4.22 14.24 4.22 14.24 3.66 14.56 3.66 ;
        POLYGON  8.27 4.54 5.82 4.54 5.82 4.22 7.95 4.22 7.95 1.88 8.27 1.88 ;
        POLYGON  7.56 2.92 7.48 2.92 7.48 3.90 2.58 3.90 2.58 4.54 2.26 4.54
                 2.26 1.28 2.58 1.28 2.58 3.58 7.16 3.58 7.16 2.60 7.56 2.60 ;
        POLYGON  6.70 3.26 6.30 3.26 6.30 2.94 6.38 2.94 6.38 2.62 5.26 2.62
                 5.26 2.30 6.38 2.30 6.38 1.88 6.70 1.88 ;
        POLYGON  5.78 3.26 4.38 3.26 4.38 2.62 2.90 2.62 2.90 2.30 4.38 2.30
                 4.38 1.66 5.70 1.66 5.70 1.98 4.70 1.98 4.70 2.94 5.78 2.94 ;
        RECT  3.05 1.26 4.06 1.58 ;
        RECT  2.96 4.22 4.06 4.54 ;
        POLYGON  1.88 1.94 0.18 1.94 0.18 1.44 0.50 1.44 0.50 1.62 1.56 1.62
                 1.56 1.60 1.88 1.60 ;
        POLYGON  1.88 4.54 1.56 4.54 1.56 3.76 0.50 3.76 0.50 4.48 0.18 4.48
                 0.18 3.44 1.88 3.44 ;
    END
END gclklatn_8

MACRO gclklatn_4
    CLASS CORE ;
    FOREIGN gclklatn_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.64 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.81  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.09 2.40 8.61 2.40 8.61 1.54 6.02 1.54 6.02 1.22 8.93 1.22
                 8.93 1.94 10.09 1.94 ;
        END
    END ck
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END g
    PIN gck
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.79  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  15.94 4.44 15.62 4.44 15.62 3.68 14.54 3.68 14.54 4.44
                 14.22 4.44 14.22 3.68 13.14 3.68 13.14 4.44 12.82 4.44
                 12.82 3.36 15.62 3.36 15.62 1.63 12.81 1.63 12.81 1.31
                 15.94 1.31 ;
        END
    END gck
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 0.90 1.20 0.90 1.20 1.30 0.88 1.30 0.88 0.90 0.00 0.90
                 0.00 -0.90 16.64 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.13 1.20 4.13
                 1.20 4.86 4.53 4.86 4.53 4.60 4.85 4.60 4.85 4.86 9.33 4.86
                 9.33 3.99 9.65 3.99 9.65 4.86 13.52 4.86 13.52 4.11 13.84 4.11
                 13.84 4.86 14.92 4.86 14.92 4.12 15.24 4.12 15.24 4.86
                 16.64 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  14.57 2.58 11.03 2.58 11.03 2.98 12.47 2.98 12.47 3.30
                 12.46 3.30 12.46 4.54 12.14 4.54 12.14 3.30 11.03 3.30
                 11.03 3.88 10.71 3.88 10.71 1.54 9.25 1.54 9.25 1.22
                 12.37 1.22 12.37 1.54 11.03 1.54 11.03 2.26 14.57 2.26 ;
        POLYGON  11.76 4.54 10.03 4.54 10.03 3.30 8.95 3.30 8.95 4.54 8.63 4.54
                 8.63 2.98 10.35 2.98 10.35 4.22 11.44 4.22 11.44 3.62
                 11.76 3.62 ;
        POLYGON  8.27 4.54 5.82 4.54 5.82 4.22 7.95 4.22 7.95 1.88 8.27 1.88 ;
        POLYGON  7.56 2.92 7.48 2.92 7.48 3.90 2.58 3.90 2.58 4.54 2.26 4.54
                 2.26 1.28 2.58 1.28 2.58 3.58 7.16 3.58 7.16 2.60 7.56 2.60 ;
        POLYGON  6.70 3.26 6.30 3.26 6.30 2.94 6.38 2.94 6.38 2.62 5.26 2.62
                 5.26 2.30 6.38 2.30 6.38 1.88 6.70 1.88 ;
        POLYGON  5.78 3.26 4.38 3.26 4.38 2.62 2.90 2.62 2.90 2.30 4.38 2.30
                 4.38 1.66 5.70 1.66 5.70 1.98 4.70 1.98 4.70 2.94 5.78 2.94 ;
        RECT  3.05 1.26 4.06 1.58 ;
        RECT  2.96 4.22 4.06 4.54 ;
        POLYGON  1.88 1.94 0.18 1.94 0.18 1.44 0.50 1.44 0.50 1.62 1.56 1.62
                 1.56 1.60 1.88 1.60 ;
        POLYGON  1.88 4.54 1.56 4.54 1.56 3.76 0.50 3.76 0.50 4.48 0.18 4.48
                 0.18 3.44 1.88 3.44 ;
    END
END gclklatn_4

MACRO gclklatn_2
    CLASS CORE ;
    FOREIGN gclklatn_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 13.44 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.44 2.40 8.59 2.40 8.59 1.54 6.02 1.54 6.02 1.22 8.91 1.22
                 8.91 1.94 9.44 1.94 ;
        END
    END ck
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END g
    PIN gck
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.04  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  13.15 3.80 13.14 3.80 13.14 4.44 12.82 4.44 12.82 3.68
                 11.74 3.68 11.74 4.44 11.42 4.44 11.42 3.36 12.82 3.36
                 12.82 1.63 11.41 1.63 11.41 1.31 13.15 1.31 ;
        END
    END gck
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  13.44 0.90 10.95 0.90 10.95 1.54 10.63 1.54 10.63 0.90
                 1.20 0.90 1.20 1.30 0.88 1.30 0.88 0.90 0.00 0.90 0.00 -0.90
                 13.44 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  13.44 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.13 1.20 4.13
                 1.20 4.86 4.53 4.86 4.53 4.60 4.85 4.60 4.85 4.86 8.63 4.86
                 8.63 3.32 8.95 3.32 8.95 4.86 12.12 4.86 12.12 4.11 12.44 4.11
                 12.44 4.86 13.44 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  12.44 2.58 11.06 2.58 11.06 4.54 10.74 4.54 10.74 2.58
                 10.63 2.58 9.93 1.88 9.93 1.22 10.25 1.22 10.25 1.74
                 10.77 2.26 12.44 2.26 ;
        POLYGON  10.33 4.54 9.33 4.54 9.33 3.04 9.65 3.04 9.65 4.22 10.33 4.22 ;
        POLYGON  8.27 4.54 5.82 4.54 5.82 4.22 7.95 4.22 7.95 1.88 8.27 1.88 ;
        POLYGON  7.56 2.92 7.48 2.92 7.48 3.90 2.58 3.90 2.58 4.54 2.26 4.54
                 2.26 1.28 2.58 1.28 2.58 3.58 7.16 3.58 7.16 2.60 7.56 2.60 ;
        POLYGON  6.70 3.26 6.30 3.26 6.30 2.94 6.38 2.94 6.38 2.62 5.26 2.62
                 5.26 2.30 6.38 2.30 6.38 1.88 6.70 1.88 ;
        POLYGON  5.78 3.26 4.38 3.26 4.38 2.62 2.90 2.62 2.90 2.30 4.38 2.30
                 4.38 1.66 5.70 1.66 5.70 1.98 4.70 1.98 4.70 2.94 5.78 2.94 ;
        RECT  3.05 1.26 4.06 1.58 ;
        RECT  2.96 4.22 4.06 4.54 ;
        POLYGON  1.88 1.94 0.18 1.94 0.18 1.44 0.50 1.44 0.50 1.62 1.56 1.62
                 1.56 1.60 1.88 1.60 ;
        POLYGON  1.88 4.54 1.56 4.54 1.56 3.76 0.50 3.76 0.50 4.48 0.18 4.48
                 0.18 3.44 1.88 3.44 ;
    END
END gclklatn_2

MACRO gclklatn_1
    CLASS CORE ;
    FOREIGN gclklatn_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.80 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.44 2.40 8.59 2.40 8.59 1.54 6.02 1.54 6.02 1.22 8.91 1.22
                 8.91 1.94 9.39 1.94 9.39 2.08 9.44 2.08 ;
        END
    END ck
    PIN g
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.84 3.04 ;
        END
    END g
    PIN gck
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.64 3.68 12.44 3.68 12.44 4.44 12.12 4.44 12.12 3.36
                 12.16 3.36 12.16 1.78 12.11 1.78 12.11 1.46 12.48 1.46
                 12.48 3.36 12.64 3.36 ;
        END
    END gck
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  12.80 0.90 11.73 0.90 11.73 1.78 11.41 1.78 11.41 0.90
                 10.95 0.90 10.95 1.54 10.63 1.54 10.63 0.90 1.20 0.90
                 1.20 1.30 0.88 1.30 0.88 0.90 0.00 0.90 0.00 -0.90 12.80 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  12.80 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.13 1.20 4.13
                 1.20 4.86 4.53 4.86 4.53 4.60 4.85 4.60 4.85 4.86 8.63 4.86
                 8.63 3.32 8.95 3.32 8.95 4.86 11.42 4.86 11.42 4.12 11.74 4.12
                 11.74 4.86 12.80 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  11.84 2.58 11.06 2.58 11.06 4.54 10.74 4.54 10.74 2.58
                 10.63 2.58 9.93 1.88 9.93 1.22 10.25 1.22 10.25 1.74
                 10.77 2.26 11.84 2.26 ;
        POLYGON  10.33 4.54 9.33 4.54 9.33 3.04 9.65 3.04 9.65 4.22 10.33 4.22 ;
        POLYGON  8.27 4.54 5.82 4.54 5.82 4.22 7.95 4.22 7.95 1.88 8.27 1.88 ;
        POLYGON  7.56 2.92 7.48 2.92 7.48 3.90 2.58 3.90 2.58 4.54 2.26 4.54
                 2.26 1.28 2.58 1.28 2.58 3.58 7.16 3.58 7.16 2.60 7.56 2.60 ;
        POLYGON  6.70 3.26 6.30 3.26 6.30 2.94 6.38 2.94 6.38 2.62 5.26 2.62
                 5.26 2.30 6.38 2.30 6.38 1.88 6.70 1.88 ;
        POLYGON  5.78 3.26 4.38 3.26 4.38 2.62 2.90 2.62 2.90 2.30 4.38 2.30
                 4.38 1.66 5.70 1.66 5.70 1.98 4.70 1.98 4.70 2.94 5.78 2.94 ;
        RECT  3.05 1.26 4.06 1.58 ;
        RECT  2.96 4.22 4.06 4.54 ;
        POLYGON  1.88 1.94 0.18 1.94 0.18 1.44 0.50 1.44 0.50 1.62 1.56 1.62
                 1.56 1.60 1.88 1.60 ;
        POLYGON  1.88 4.54 1.56 4.54 1.56 3.76 0.50 3.76 0.50 4.48 0.18 4.48
                 0.18 3.44 1.88 3.44 ;
    END
END gclklatn_1

MACRO fill_8
    CLASS CORE SPACER ;
    FOREIGN fill_8 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 0.90 4.70 0.90 4.70 1.30 4.38 1.30 4.38 0.90 0.74 0.90
                 0.74 1.30 0.42 1.30 0.42 0.90 0.00 0.90 0.00 -0.90 5.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 6.66 0.00 6.66 0.00 4.86 0.42 4.86 0.42 3.34 0.74 3.34
                 0.74 4.86 4.38 4.86 4.38 3.34 4.70 3.34 4.70 4.86 5.12 4.86 ;
        END
    END vdd!
END fill_8

MACRO fill_4
    CLASS CORE SPACER ;
    FOREIGN fill_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.56 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  2.56 0.90 2.14 0.90 2.14 1.30 1.82 1.30 1.82 0.90 0.74 0.90
                 0.74 1.30 0.42 1.30 0.42 0.90 0.00 0.90 0.00 -0.90 2.56 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  2.56 6.66 0.00 6.66 0.00 4.86 0.42 4.86 0.42 3.34 0.74 3.34
                 0.74 4.86 1.82 4.86 1.82 3.34 2.14 3.34 2.14 4.86 2.56 4.86 ;
        END
    END vdd!
END fill_4

MACRO fill_32
    CLASS CORE SPACER ;
    FOREIGN fill_32 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 20.48 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 0.90 20.06 0.90 20.06 1.30 19.74 1.30 19.74 0.90
                 0.74 0.90 0.74 1.30 0.42 1.30 0.42 0.90 0.00 0.90 0.00 -0.90
                 20.48 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 6.66 0.00 6.66 0.00 4.86 0.42 4.86 0.42 3.34 0.74 3.34
                 0.74 4.86 19.74 4.86 19.74 3.34 20.06 3.34 20.06 4.86
                 20.48 4.86 ;
        END
    END vdd!
END fill_32

MACRO fill_2
    CLASS CORE SPACER ;
    FOREIGN fill_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 1.28 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 1.28 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 1.28 6.66 ;
        END
    END vdd!
END fill_2

MACRO fill_16
    CLASS CORE SPACER ;
    FOREIGN fill_16 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.24 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  10.24 0.90 9.82 0.90 9.82 1.30 9.50 1.30 9.50 0.90 0.74 0.90
                 0.74 1.30 0.42 1.30 0.42 0.90 0.00 0.90 0.00 -0.90 10.24 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  10.24 6.66 0.00 6.66 0.00 4.86 0.42 4.86 0.42 3.34 0.74 3.34
                 0.74 4.86 9.50 4.86 9.50 3.34 9.82 3.34 9.82 4.86 10.24 4.86 ;
        END
    END vdd!
END fill_16

MACRO fill_1
    CLASS CORE SPACER ;
    FOREIGN fill_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 0.64 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 0.64 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 0.64 6.66 ;
        END
    END vdd!
END fill_1

MACRO exor4_4
    CLASS CORE ;
    FOREIGN exor4_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  19.84 2.58 20.32 3.22 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  18.56 2.72 19.10 3.22 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.86 2.72 2.40 3.22 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.58 1.12 3.22 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.56 1.88 14.02 1.88 14.02 4.54 13.69 4.54 13.69 3.68
                 12.63 3.68 12.63 4.54 12.30 4.54 12.30 3.36 13.69 3.36
                 13.69 1.88 12.84 1.88 12.84 1.22 13.16 1.22 13.16 1.56
                 14.24 1.56 14.24 1.22 14.56 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 0.90 18.70 0.90 18.70 1.54 18.38 1.54 18.38 0.90
                 13.86 0.90 13.86 1.22 13.54 1.22 13.54 0.90 8.88 0.90
                 8.88 1.18 8.56 1.18 8.56 0.90 2.58 0.90 2.58 1.54 2.26 1.54
                 2.26 0.90 0.00 0.90 0.00 -0.90 21.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.62 1.32 4.62
                 1.32 4.86 7.30 4.86 7.30 4.62 7.62 4.62 7.62 4.86 10.86 4.86
                 10.86 4.62 11.18 4.62 11.18 4.86 13.00 4.86 13.00 4.61
                 13.32 4.61 13.32 4.86 19.64 4.86 19.64 4.61 19.96 4.61
                 19.96 4.86 21.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.96 4.23 18.94 4.23 18.94 3.91 20.64 3.91 20.64 2.18
                 16.16 2.18 16.16 2.50 15.84 2.50 15.84 1.86 20.64 1.86
                 20.64 1.54 20.46 1.54 20.46 1.22 20.96 1.22 ;
        RECT  19.08 1.22 20.08 1.54 ;
        POLYGON  18.58 4.54 14.35 4.54 14.35 4.22 14.92 4.22 14.92 1.22
                 15.24 1.22 15.24 4.22 18.26 4.22 18.26 3.58 18.58 3.58 ;
        RECT  15.62 1.22 18.02 1.54 ;
        RECT  16.80 2.94 17.88 3.90 ;
        POLYGON  13.16 2.52 12.48 2.52 12.48 2.90 11.94 2.90 11.94 4.27
                 8.68 4.27 8.68 2.94 9.00 2.94 9.00 3.95 11.62 3.95 11.62 2.58
                 12.16 2.58 12.16 1.22 12.48 1.22 12.48 2.20 13.16 2.20 ;
        POLYGON  11.84 2.26 11.52 2.26 11.52 2.18 8.32 2.18 8.32 4.30 6.60 4.30
                 6.60 3.98 8.00 3.98 8.00 2.18 6.48 2.18 6.48 1.22 6.80 1.22
                 6.80 1.86 11.84 1.86 ;
        RECT  9.30 1.22 11.78 1.54 ;
        POLYGON  10.43 3.60 9.38 3.60 9.38 3.28 10.10 3.28 10.10 2.64
                 10.43 2.64 ;
        RECT  7.18 1.22 8.18 1.54 ;
        POLYGON  7.04 3.22 6.12 3.22 6.12 4.54 2.38 4.54 2.38 3.58 2.70 3.58
                 2.70 4.22 5.80 4.22 5.80 1.22 6.12 1.22 6.12 2.90 7.04 2.90 ;
        RECT  2.94 1.22 5.42 1.54 ;
        POLYGON  5.20 2.50 4.88 2.50 4.88 2.18 0.48 2.18 0.48 3.98 2.02 3.98
                 2.02 4.30 0.16 4.30 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 1.86 5.20 1.86 ;
        RECT  3.08 2.94 4.24 3.90 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END exor4_4

MACRO exor4_2
    CLASS CORE ;
    FOREIGN exor4_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 20.48 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  19.18 2.58 19.68 3.22 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  17.86 2.72 18.40 3.22 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.86 2.72 2.40 3.22 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.58 1.12 3.22 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  13.86 3.68 13.32 3.68 13.32 4.54 12.96 4.54 12.96 3.36
                 13.54 3.36 13.54 1.22 13.86 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 0.90 18.00 0.90 18.00 1.54 17.68 1.54 17.68 0.90
                 13.16 0.90 13.16 1.22 12.84 1.22 12.84 0.90 8.88 0.90
                 8.88 1.18 8.56 1.18 8.56 0.90 2.58 0.90 2.58 1.54 2.26 1.54
                 2.26 0.90 0.00 0.90 0.00 -0.90 20.48 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.62 1.32 4.62
                 1.32 4.86 7.30 4.86 7.30 4.62 7.62 4.62 7.62 4.86 10.86 4.86
                 10.86 4.62 11.18 4.62 11.18 4.86 12.30 4.86 12.30 4.61
                 12.62 4.61 12.62 4.86 18.94 4.86 18.94 4.61 19.26 4.61
                 19.26 4.86 20.48 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.32 4.23 18.24 4.23 18.24 3.91 20.00 3.91 20.00 2.18
                 15.46 2.18 15.46 2.50 15.14 2.50 15.14 1.86 20.00 1.86
                 20.00 1.54 19.76 1.54 19.76 1.22 20.32 1.22 ;
        RECT  18.38 1.22 19.38 1.54 ;
        POLYGON  17.88 4.54 13.65 4.54 13.65 4.22 14.22 4.22 14.22 1.22
                 14.54 1.22 14.54 4.22 17.56 4.22 17.56 3.58 17.88 3.58 ;
        RECT  14.92 1.22 17.32 1.54 ;
        RECT  16.10 2.94 17.18 3.90 ;
        POLYGON  13.20 2.52 12.48 2.52 12.48 2.90 11.94 2.90 11.94 4.27
                 8.68 4.27 8.68 2.94 9.00 2.94 9.00 3.95 11.62 3.95 11.62 2.58
                 12.16 2.58 12.16 1.22 12.48 1.22 12.48 2.20 13.20 2.20 ;
        POLYGON  11.84 2.26 11.52 2.26 11.52 2.18 8.32 2.18 8.32 4.30 6.60 4.30
                 6.60 3.98 8.00 3.98 8.00 2.18 6.48 2.18 6.48 1.22 6.80 1.22
                 6.80 1.86 11.84 1.86 ;
        RECT  9.30 1.22 11.78 1.54 ;
        POLYGON  10.43 3.60 9.38 3.60 9.38 3.28 10.10 3.28 10.10 2.64
                 10.43 2.64 ;
        RECT  7.18 1.22 8.18 1.54 ;
        POLYGON  7.04 3.22 6.12 3.22 6.12 4.54 2.38 4.54 2.38 3.58 2.70 3.58
                 2.70 4.22 5.80 4.22 5.80 1.22 6.12 1.22 6.12 2.90 7.04 2.90 ;
        RECT  2.94 1.22 5.42 1.54 ;
        POLYGON  5.20 2.50 4.88 2.50 4.88 2.18 0.48 2.18 0.48 3.98 2.02 3.98
                 2.02 4.30 0.16 4.30 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 1.86 5.20 1.86 ;
        RECT  3.08 2.94 4.24 3.90 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END exor4_2

MACRO exor4_1
    CLASS CORE ;
    FOREIGN exor4_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 20.48 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  19.18 2.58 19.68 3.22 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  17.86 2.72 18.40 3.22 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.86 2.72 2.40 3.22 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.58 1.12 3.22 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  13.86 3.68 13.32 3.68 13.32 4.54 12.96 4.54 12.96 3.36
                 13.54 3.36 13.54 1.22 13.86 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 0.90 18.00 0.90 18.00 1.54 17.68 1.54 17.68 0.90
                 13.16 0.90 13.16 1.27 12.84 1.27 12.84 0.90 8.88 0.90
                 8.88 1.18 8.56 1.18 8.56 0.90 2.58 0.90 2.58 1.54 2.26 1.54
                 2.26 0.90 0.00 0.90 0.00 -0.90 20.48 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.62 1.32 4.62
                 1.32 4.86 7.30 4.86 7.30 4.62 7.62 4.62 7.62 4.86 10.86 4.86
                 10.86 4.62 11.18 4.62 11.18 4.86 12.30 4.86 12.30 4.61
                 12.62 4.61 12.62 4.86 18.94 4.86 18.94 4.61 19.26 4.61
                 19.26 4.86 20.48 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.32 4.23 18.24 4.23 18.24 3.91 20.00 3.91 20.00 2.18
                 15.46 2.18 15.46 2.50 15.14 2.50 15.14 1.86 20.00 1.86
                 20.00 1.54 19.76 1.54 19.76 1.22 20.32 1.22 ;
        RECT  18.38 1.22 19.38 1.54 ;
        POLYGON  17.88 4.54 13.65 4.54 13.65 4.22 14.22 4.22 14.22 1.22
                 14.54 1.22 14.54 4.22 17.56 4.22 17.56 3.58 17.88 3.58 ;
        RECT  14.92 1.22 17.32 1.54 ;
        RECT  16.10 2.94 17.18 3.90 ;
        POLYGON  13.20 2.52 12.48 2.52 12.48 2.90 11.94 2.90 11.94 4.27
                 8.68 4.27 8.68 2.94 9.00 2.94 9.00 3.95 11.62 3.95 11.62 2.58
                 12.16 2.58 12.16 1.22 12.48 1.22 12.48 2.20 13.20 2.20 ;
        POLYGON  11.84 2.26 11.52 2.26 11.52 2.18 8.32 2.18 8.32 4.30 6.60 4.30
                 6.60 3.98 8.00 3.98 8.00 2.18 6.48 2.18 6.48 1.22 6.80 1.22
                 6.80 1.86 11.84 1.86 ;
        RECT  9.30 1.22 11.78 1.54 ;
        POLYGON  10.43 3.60 9.38 3.60 9.38 3.28 10.10 3.28 10.10 2.64
                 10.43 2.64 ;
        RECT  7.18 1.22 8.18 1.54 ;
        POLYGON  7.04 3.22 6.12 3.22 6.12 4.54 2.38 4.54 2.38 3.58 2.70 3.58
                 2.70 4.22 5.80 4.22 5.80 1.22 6.12 1.22 6.12 2.90 7.04 2.90 ;
        RECT  2.94 1.22 5.42 1.54 ;
        POLYGON  5.20 2.50 4.88 2.50 4.88 2.18 0.48 2.18 0.48 3.98 2.02 3.98
                 2.02 4.30 0.16 4.30 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 1.86 5.20 1.86 ;
        RECT  3.08 2.94 4.24 3.90 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END exor4_1

MACRO exor3_4
    CLASS CORE ;
    FOREIGN exor3_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.64 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  11.40 2.72 12.04 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.58 1.12 3.22 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.86 2.72 2.40 3.22 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  15.88 4.54 15.56 4.54 15.56 3.82 14.48 3.82 14.48 4.54
                 14.16 4.54 14.16 3.50 15.56 3.50 15.56 3.04 15.52 3.04
                 15.52 2.72 15.56 2.72 15.56 2.17 14.16 2.17 14.16 1.22
                 14.48 1.22 14.48 1.85 15.56 1.85 15.56 1.22 15.88 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 0.90 15.18 0.90 15.18 1.48 14.86 1.48 14.86 0.90
                 10.26 0.90 10.26 1.54 9.94 1.54 9.94 0.90 6.80 0.90 6.80 1.54
                 6.48 1.54 6.48 0.90 2.58 0.90 2.58 1.54 2.26 1.54 2.26 0.90
                 0.00 0.90 0.00 -0.90 16.64 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.62 1.32 4.62
                 1.32 4.86 6.48 4.86 6.48 4.22 6.80 4.22 6.80 4.86 8.68 4.86
                 8.68 4.62 9.00 4.62 9.00 4.86 14.86 4.86 14.86 4.21 15.18 4.21
                 15.18 4.86 16.64 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  15.14 2.98 13.80 2.98 13.80 4.54 10.06 4.54 10.06 2.94
                 10.38 2.94 10.38 4.22 13.48 4.22 13.48 1.22 13.80 1.22
                 13.80 2.66 15.14 2.66 ;
        POLYGON  13.16 2.50 12.84 2.50 12.84 2.18 9.70 2.18 9.70 4.54 9.38 4.54
                 9.38 4.30 8.30 4.30 8.30 4.54 7.98 4.54 7.98 3.58 8.30 3.58
                 8.30 3.98 9.38 3.98 9.38 2.18 7.86 2.18 7.86 1.22 8.18 1.22
                 8.18 1.86 13.16 1.86 ;
        RECT  10.62 1.22 13.10 1.54 ;
        POLYGON  12.30 3.90 10.76 3.90 10.76 2.94 11.08 2.94 11.08 3.58
                 12.30 3.58 ;
        RECT  8.56 1.22 9.56 1.54 ;
        POLYGON  8.42 3.22 7.50 3.22 7.50 4.54 7.18 4.54 7.18 1.22 7.50 1.22
                 7.50 2.90 8.42 2.90 ;
        POLYGON  6.86 2.92 6.12 2.92 6.12 4.54 2.38 4.54 2.38 3.58 2.70 3.58
                 2.70 4.22 5.80 4.22 5.80 1.22 6.12 1.22 6.12 2.60 6.86 2.60 ;
        RECT  2.94 1.22 5.42 1.54 ;
        POLYGON  5.20 2.50 4.88 2.50 4.88 2.18 0.48 2.18 0.48 3.58 0.50 3.58
                 0.50 3.98 1.70 3.98 1.70 3.58 2.02 3.58 2.02 4.54 1.70 4.54
                 1.70 4.30 0.50 4.30 0.50 4.54 0.18 4.54 0.18 4.30 0.16 4.30
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 1.86 5.20 1.86 ;
        RECT  3.08 2.94 4.24 3.90 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END exor3_4

MACRO exor3_2
    CLASS CORE ;
    FOREIGN exor3_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.36 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  11.40 2.72 12.04 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.58 1.12 3.22 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.86 2.72 2.40 3.22 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  15.20 3.04 15.18 3.04 15.18 4.54 14.86 4.54 14.86 1.22
                 15.18 1.22 15.18 2.72 15.20 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  15.36 0.90 14.48 0.90 14.48 1.54 14.16 1.54 14.16 0.90
                 10.26 0.90 10.26 1.54 9.94 1.54 9.94 0.90 6.80 0.90 6.80 1.54
                 6.48 1.54 6.48 0.90 2.58 0.90 2.58 1.54 2.26 1.54 2.26 0.90
                 0.00 0.90 0.00 -0.90 15.36 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  15.36 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.62 1.32 4.62
                 1.32 4.86 6.48 4.86 6.48 4.22 6.80 4.22 6.80 4.86 8.68 4.86
                 8.68 4.62 9.00 4.62 9.00 4.86 14.16 4.86 14.16 3.58 14.48 3.58
                 14.48 4.86 15.36 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  14.54 2.98 13.80 2.98 13.80 4.54 10.06 4.54 10.06 2.94
                 10.38 2.94 10.38 4.22 13.48 4.22 13.48 1.22 13.80 1.22
                 13.80 2.66 14.54 2.66 ;
        POLYGON  13.16 2.50 12.84 2.50 12.84 2.18 9.70 2.18 9.70 4.54 9.38 4.54
                 9.38 4.30 8.30 4.30 8.30 4.54 7.98 4.54 7.98 3.58 8.30 3.58
                 8.30 3.98 9.38 3.98 9.38 2.18 7.86 2.18 7.86 1.22 8.18 1.22
                 8.18 1.86 13.16 1.86 ;
        RECT  10.62 1.22 13.10 1.54 ;
        POLYGON  12.30 3.90 10.76 3.90 10.76 2.94 11.08 2.94 11.08 3.58
                 12.30 3.58 ;
        RECT  8.56 1.22 9.56 1.54 ;
        POLYGON  8.42 3.22 7.50 3.22 7.50 4.54 7.18 4.54 7.18 1.22 7.50 1.22
                 7.50 2.90 8.42 2.90 ;
        POLYGON  6.86 2.92 6.12 2.92 6.12 4.54 2.38 4.54 2.38 3.58 2.70 3.58
                 2.70 4.22 5.80 4.22 5.80 1.22 6.12 1.22 6.12 2.60 6.86 2.60 ;
        RECT  2.94 1.22 5.42 1.54 ;
        POLYGON  5.20 2.50 4.88 2.50 4.88 2.18 0.48 2.18 0.48 3.58 0.50 3.58
                 0.50 3.98 1.70 3.98 1.70 3.58 2.02 3.58 2.02 4.54 1.70 4.54
                 1.70 4.30 0.50 4.30 0.50 4.54 0.18 4.54 0.18 4.30 0.16 4.30
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 1.86 5.20 1.86 ;
        RECT  3.08 2.94 4.24 3.90 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END exor3_2

MACRO exor3_1
    CLASS CORE ;
    FOREIGN exor3_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.36 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  11.40 2.72 12.04 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.58 1.12 3.22 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.86 2.72 2.40 3.22 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  15.20 3.04 15.18 3.04 15.18 4.54 14.86 4.54 14.86 1.22
                 15.18 1.22 15.18 2.72 15.20 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  15.36 0.90 14.48 0.90 14.48 1.54 14.16 1.54 14.16 0.90
                 10.26 0.90 10.26 1.54 9.94 1.54 9.94 0.90 6.80 0.90 6.80 1.54
                 6.48 1.54 6.48 0.90 2.58 0.90 2.58 1.54 2.26 1.54 2.26 0.90
                 0.00 0.90 0.00 -0.90 15.36 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  15.36 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.62 1.32 4.62
                 1.32 4.86 6.48 4.86 6.48 4.22 6.80 4.22 6.80 4.86 8.68 4.86
                 8.68 4.62 9.00 4.62 9.00 4.86 14.16 4.86 14.16 4.22 14.48 4.22
                 14.48 4.86 15.36 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  14.54 2.92 13.80 2.92 13.80 4.54 10.06 4.54 10.06 2.94
                 10.38 2.94 10.38 4.22 13.48 4.22 13.48 1.22 13.80 1.22
                 13.80 2.60 14.54 2.60 ;
        POLYGON  13.16 2.50 12.84 2.50 12.84 2.18 9.70 2.18 9.70 4.30 7.98 4.30
                 7.98 3.98 9.38 3.98 9.38 2.18 7.86 2.18 7.86 1.22 8.18 1.22
                 8.18 1.86 13.16 1.86 ;
        RECT  10.62 1.22 13.10 1.54 ;
        POLYGON  12.30 3.90 10.76 3.90 10.76 2.94 11.08 2.94 11.08 3.58
                 12.30 3.58 ;
        RECT  8.56 1.22 9.56 1.54 ;
        POLYGON  8.42 3.22 7.50 3.22 7.50 4.54 7.18 4.54 7.18 1.22 7.50 1.22
                 7.50 2.90 8.42 2.90 ;
        POLYGON  6.86 2.92 6.12 2.92 6.12 4.54 2.38 4.54 2.38 3.58 2.70 3.58
                 2.70 4.22 5.80 4.22 5.80 1.22 6.12 1.22 6.12 2.60 6.86 2.60 ;
        RECT  2.94 1.22 5.42 1.54 ;
        POLYGON  5.20 2.50 4.88 2.50 4.88 2.18 0.48 2.18 0.48 3.98 2.02 3.98
                 2.02 4.30 0.16 4.30 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 1.86 5.20 1.86 ;
        RECT  3.08 2.94 4.24 3.90 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END exor3_1

MACRO exor2_4
    CLASS CORE ;
    FOREIGN exor2_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.96 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.58 1.12 3.22 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.86 2.72 2.40 3.22 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.20 4.54 7.88 4.54 7.88 3.78 6.80 3.78 6.80 4.54 6.48 4.54
                 6.48 3.46 7.88 3.46 7.88 3.04 7.84 3.04 7.84 2.72 7.88 2.72
                 7.88 2.14 6.48 2.14 6.48 1.22 6.80 1.22 6.80 1.82 7.88 1.82
                 7.88 1.22 8.20 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.96 0.90 7.50 0.90 7.50 1.46 7.18 1.46 7.18 0.90 2.58 0.90
                 2.58 1.54 2.26 1.54 2.26 0.90 0.00 0.90 0.00 -0.90 8.96 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  8.96 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.62 1.32 4.62
                 1.32 4.86 7.18 4.86 7.18 4.21 7.50 4.21 7.50 4.86 8.96 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  7.40 2.98 6.12 2.98 6.12 4.54 2.38 4.54 2.38 3.58 2.70 3.58
                 2.70 4.22 5.80 4.22 5.80 1.22 6.12 1.22 6.12 2.66 7.40 2.66 ;
        RECT  2.94 1.22 5.42 1.54 ;
        POLYGON  5.20 2.50 4.88 2.50 4.88 2.18 0.48 2.18 0.48 3.98 2.02 3.98
                 2.02 4.30 0.16 4.30 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 1.86 5.20 1.86 ;
        RECT  3.08 2.94 4.08 3.90 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END exor2_4

MACRO exor2_2
    CLASS CORE ;
    FOREIGN exor2_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.58 1.12 3.22 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.86 2.72 2.40 3.22 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.52 3.04 7.50 3.04 7.50 4.54 7.18 4.54 7.18 1.22 7.50 1.22
                 7.50 2.72 7.52 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 0.90 6.80 0.90 6.80 1.54 6.48 1.54 6.48 0.90 2.58 0.90
                 2.58 1.54 2.26 1.54 2.26 0.90 0.00 0.90 0.00 -0.90 7.68 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.62 1.32 4.62
                 1.32 4.86 6.48 4.86 6.48 3.58 6.80 3.58 6.80 4.86 7.68 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  6.86 2.98 6.12 2.98 6.12 4.54 2.38 4.54 2.38 3.58 2.70 3.58
                 2.70 4.22 5.80 4.22 5.80 1.22 6.12 1.22 6.12 2.66 6.86 2.66 ;
        RECT  2.94 1.22 5.42 1.54 ;
        POLYGON  5.20 2.50 4.88 2.50 4.88 2.18 0.48 2.18 0.48 3.98 2.02 3.98
                 2.02 4.30 0.16 4.30 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 1.86 5.20 1.86 ;
        RECT  3.08 2.94 4.08 3.90 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END exor2_2

MACRO exor2_1
    CLASS CORE ;
    FOREIGN exor2_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.58 1.12 3.22 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.86 2.72 2.40 3.22 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.52 3.04 7.50 3.04 7.50 4.54 7.18 4.54 7.18 1.22 7.50 1.22
                 7.50 2.72 7.52 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 0.90 6.80 0.90 6.80 1.54 6.48 1.54 6.48 0.90 2.58 0.90
                 2.58 1.54 2.26 1.54 2.26 0.90 0.00 0.90 0.00 -0.90 7.68 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.62 1.32 4.62
                 1.32 4.86 6.48 4.86 6.48 4.34 6.80 4.34 6.80 4.86 7.68 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  6.86 2.92 6.12 2.92 6.12 4.54 2.38 4.54 2.38 3.58 2.70 3.58
                 2.70 4.22 5.80 4.22 5.80 1.22 6.12 1.22 6.12 2.60 6.86 2.60 ;
        RECT  2.94 1.22 5.42 1.54 ;
        POLYGON  5.20 2.50 4.88 2.50 4.88 2.18 0.48 2.18 0.48 3.98 2.02 3.98
                 2.02 4.30 0.16 4.30 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 1.86 5.20 1.86 ;
        RECT  3.08 2.94 4.08 3.90 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END exor2_1

MACRO exnor4_4
    CLASS CORE ;
    FOREIGN exnor4_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  21.22 2.58 21.60 3.22 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  19.94 2.72 20.48 3.22 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.86 2.72 2.40 3.22 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.58 1.12 3.22 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  15.94 1.88 15.40 1.88 15.40 4.54 15.07 4.54 15.07 3.68
                 14.56 3.68 14.56 3.92 14.01 3.92 14.01 4.54 13.68 4.54
                 13.68 3.60 14.24 3.60 14.24 3.36 15.07 3.36 15.07 1.88
                 14.22 1.88 14.22 1.22 14.54 1.22 14.54 1.56 15.62 1.56
                 15.62 1.22 15.94 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  22.40 0.90 20.08 0.90 20.08 1.54 19.76 1.54 19.76 0.90
                 15.24 0.90 15.24 1.22 14.92 1.22 14.92 0.90 13.86 0.90
                 13.86 1.16 13.54 1.16 13.54 0.90 8.88 0.90 8.88 1.18 8.56 1.18
                 8.56 0.90 2.58 0.90 2.58 1.54 2.26 1.54 2.26 0.90 0.00 0.90
                 0.00 -0.90 22.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  22.40 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.62 1.32 4.62
                 1.32 4.86 7.30 4.86 7.30 4.62 7.62 4.62 7.62 4.86 10.86 4.86
                 10.86 4.62 11.18 4.62 11.18 4.86 13.00 4.86 13.00 4.60
                 13.32 4.60 13.32 4.86 14.38 4.86 14.38 4.61 14.70 4.61
                 14.70 4.86 21.02 4.86 21.02 4.61 21.34 4.61 21.34 4.86
                 22.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  22.24 4.23 20.32 4.23 20.32 3.91 21.92 3.91 21.92 2.18
                 17.54 2.18 17.54 2.50 17.22 2.50 17.22 1.86 21.92 1.86
                 21.92 1.54 21.84 1.54 21.84 1.22 22.24 1.22 ;
        RECT  20.46 1.22 21.46 1.54 ;
        POLYGON  19.96 4.54 15.73 4.54 15.73 4.22 16.30 4.22 16.30 1.22
                 16.62 1.22 16.62 4.22 19.64 4.22 19.64 3.58 19.96 3.58 ;
        RECT  17.00 1.22 19.40 1.54 ;
        RECT  18.18 2.94 19.26 3.90 ;
        POLYGON  14.74 2.52 13.68 2.52 13.68 3.25 13.36 3.25 13.36 3.92
                 12.63 3.92 12.63 4.54 12.30 4.54 12.30 3.60 13.04 3.60
                 13.04 2.93 13.36 2.93 13.36 1.88 12.84 1.88 12.84 1.22
                 13.16 1.22 13.16 1.56 13.68 1.56 13.68 2.20 14.74 2.20 ;
        POLYGON  13.03 2.52 12.48 2.52 12.48 2.90 11.94 2.90 11.94 4.27
                 8.68 4.27 8.68 2.94 9.00 2.94 9.00 3.95 11.62 3.95 11.62 2.58
                 12.16 2.58 12.16 1.22 12.48 1.22 12.48 2.20 13.03 2.20 ;
        POLYGON  11.84 2.26 11.52 2.26 11.52 2.18 8.32 2.18 8.32 4.30 6.60 4.30
                 6.60 3.98 8.00 3.98 8.00 2.18 6.48 2.18 6.48 1.22 6.80 1.22
                 6.80 1.86 11.84 1.86 ;
        RECT  9.30 1.22 11.78 1.54 ;
        POLYGON  10.43 3.60 9.38 3.60 9.38 3.28 10.10 3.28 10.10 2.64
                 10.43 2.64 ;
        RECT  7.18 1.22 8.18 1.54 ;
        POLYGON  7.04 3.22 6.12 3.22 6.12 4.54 2.38 4.54 2.38 3.58 2.70 3.58
                 2.70 4.22 5.80 4.22 5.80 1.22 6.12 1.22 6.12 2.90 7.04 2.90 ;
        RECT  2.94 1.22 5.42 1.54 ;
        POLYGON  5.20 2.50 4.88 2.50 4.88 2.18 0.48 2.18 0.48 3.98 2.02 3.98
                 2.02 4.30 0.16 4.30 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 1.86 5.20 1.86 ;
        RECT  3.08 2.94 4.24 3.90 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END exnor4_4

MACRO exnor4_2
    CLASS CORE ;
    FOREIGN exnor4_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.76 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  20.58 2.58 20.96 3.22 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  19.26 2.72 19.80 3.22 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.86 2.72 2.40 3.22 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.58 1.12 3.22 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  15.26 3.68 14.72 3.68 14.72 4.54 14.39 4.54 14.39 3.36
                 14.94 3.36 14.94 1.22 15.26 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.76 0.90 19.40 0.90 19.40 1.54 19.08 1.54 19.08 0.90
                 14.56 0.90 14.56 1.22 14.24 1.22 14.24 0.90 8.88 0.90
                 8.88 1.18 8.56 1.18 8.56 0.90 2.58 0.90 2.58 1.54 2.26 1.54
                 2.26 0.90 0.00 0.90 0.00 -0.90 21.76 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.76 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.62 1.32 4.62
                 1.32 4.86 7.30 4.86 7.30 4.62 7.62 4.62 7.62 4.86 10.86 4.86
                 10.86 4.62 11.18 4.62 11.18 4.86 12.30 4.86 12.30 4.60
                 12.62 4.60 12.62 4.86 13.70 4.86 13.70 4.61 14.02 4.61
                 14.02 4.86 20.34 4.86 20.34 4.61 20.66 4.61 20.66 4.86
                 21.76 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  21.60 4.23 19.64 4.23 19.64 3.91 21.28 3.91 21.28 2.18
                 16.86 2.18 16.86 2.50 16.54 2.50 16.54 1.86 21.28 1.86
                 21.28 1.54 21.16 1.54 21.16 1.22 21.60 1.22 ;
        RECT  19.78 1.22 20.78 1.54 ;
        POLYGON  19.28 4.54 15.05 4.54 15.05 4.22 15.62 4.22 15.62 1.22
                 15.94 1.22 15.94 4.22 18.96 4.22 18.96 3.58 19.28 3.58 ;
        RECT  16.32 1.22 18.72 1.54 ;
        RECT  17.50 2.94 18.58 3.90 ;
        POLYGON  14.60 2.52 13.68 2.52 13.68 3.25 13.36 3.25 13.36 3.92
                 13.33 3.92 13.33 4.54 13.00 4.54 13.00 3.60 13.04 3.60
                 13.04 2.93 13.36 2.93 13.36 1.54 12.84 1.54 12.84 1.22
                 13.68 1.22 13.68 2.20 14.60 2.20 ;
        POLYGON  13.03 2.52 12.48 2.52 12.48 2.90 11.94 2.90 11.94 4.27
                 8.68 4.27 8.68 2.94 9.00 2.94 9.00 3.95 11.62 3.95 11.62 2.58
                 12.16 2.58 12.16 1.22 12.48 1.22 12.48 2.20 13.03 2.20 ;
        POLYGON  11.84 2.26 11.52 2.26 11.52 2.18 8.32 2.18 8.32 4.30 6.60 4.30
                 6.60 3.98 8.00 3.98 8.00 2.18 6.48 2.18 6.48 1.22 6.80 1.22
                 6.80 1.86 11.84 1.86 ;
        RECT  9.30 1.22 11.78 1.54 ;
        POLYGON  10.43 3.60 9.38 3.60 9.38 3.28 10.10 3.28 10.10 2.64
                 10.43 2.64 ;
        RECT  7.18 1.22 8.18 1.54 ;
        POLYGON  7.04 3.22 6.12 3.22 6.12 4.54 2.38 4.54 2.38 3.58 2.70 3.58
                 2.70 4.22 5.80 4.22 5.80 1.22 6.12 1.22 6.12 2.90 7.04 2.90 ;
        RECT  2.94 1.22 5.42 1.54 ;
        POLYGON  5.20 2.50 4.88 2.50 4.88 2.18 0.48 2.18 0.48 3.98 2.02 3.98
                 2.02 4.30 0.16 4.30 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 1.86 5.20 1.86 ;
        RECT  3.08 2.94 4.24 3.90 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END exnor4_2

MACRO exnor4_1
    CLASS CORE ;
    FOREIGN exnor4_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.76 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  20.58 2.58 20.96 3.22 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  19.26 2.72 19.80 3.22 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.86 2.72 2.40 3.22 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.58 1.12 3.22 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  15.26 3.68 14.72 3.68 14.72 4.54 14.39 4.54 14.39 3.36
                 14.94 3.36 14.94 1.22 15.26 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.76 0.90 19.40 0.90 19.40 1.54 19.08 1.54 19.08 0.90
                 14.56 0.90 14.56 1.22 14.24 1.22 14.24 0.90 8.88 0.90
                 8.88 1.18 8.56 1.18 8.56 0.90 2.58 0.90 2.58 1.54 2.26 1.54
                 2.26 0.90 0.00 0.90 0.00 -0.90 21.76 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.76 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.62 1.32 4.62
                 1.32 4.86 7.30 4.86 7.30 4.62 7.62 4.62 7.62 4.86 10.86 4.86
                 10.86 4.62 11.18 4.62 11.18 4.86 12.30 4.86 12.30 4.60
                 12.62 4.60 12.62 4.86 13.70 4.86 13.70 3.99 14.02 3.99
                 14.02 4.86 20.34 4.86 20.34 4.61 20.66 4.61 20.66 4.86
                 21.76 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  21.60 4.23 19.64 4.23 19.64 3.91 21.28 3.91 21.28 2.18
                 16.86 2.18 16.86 2.50 16.54 2.50 16.54 1.86 21.28 1.86
                 21.28 1.54 21.16 1.54 21.16 1.22 21.60 1.22 ;
        RECT  19.78 1.22 20.78 1.54 ;
        POLYGON  19.28 4.54 15.05 4.54 15.05 4.22 15.62 4.22 15.62 1.22
                 15.94 1.22 15.94 4.22 18.96 4.22 18.96 3.58 19.28 3.58 ;
        RECT  16.32 1.22 18.72 1.54 ;
        RECT  17.50 2.94 18.58 3.90 ;
        POLYGON  14.60 2.52 13.68 2.52 13.68 3.25 13.36 3.25 13.36 3.92
                 13.33 3.92 13.33 4.54 13.00 4.54 13.00 3.60 13.04 3.60
                 13.04 2.93 13.36 2.93 13.36 1.54 12.84 1.54 12.84 1.22
                 13.68 1.22 13.68 2.20 14.60 2.20 ;
        POLYGON  13.03 2.52 12.48 2.52 12.48 2.90 11.94 2.90 11.94 4.27
                 8.68 4.27 8.68 2.94 9.00 2.94 9.00 3.95 11.62 3.95 11.62 2.58
                 12.16 2.58 12.16 1.22 12.48 1.22 12.48 2.20 13.03 2.20 ;
        POLYGON  11.84 2.26 11.52 2.26 11.52 2.18 8.32 2.18 8.32 4.30 6.60 4.30
                 6.60 3.98 8.00 3.98 8.00 2.18 6.48 2.18 6.48 1.22 6.80 1.22
                 6.80 1.86 11.84 1.86 ;
        RECT  9.30 1.22 11.78 1.54 ;
        POLYGON  10.43 3.60 9.38 3.60 9.38 3.28 10.10 3.28 10.10 2.64
                 10.43 2.64 ;
        RECT  7.18 1.22 8.18 1.54 ;
        POLYGON  7.04 3.22 6.12 3.22 6.12 4.54 2.38 4.54 2.38 3.58 2.70 3.58
                 2.70 4.22 5.80 4.22 5.80 1.22 6.12 1.22 6.12 2.90 7.04 2.90 ;
        RECT  2.94 1.22 5.42 1.54 ;
        POLYGON  5.20 2.50 4.88 2.50 4.88 2.18 0.48 2.18 0.48 3.98 2.02 3.98
                 2.02 4.30 0.16 4.30 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 1.86 5.20 1.86 ;
        RECT  3.08 2.94 4.24 3.90 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END exnor4_1

MACRO exnor3_4
    CLASS CORE ;
    FOREIGN exnor3_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.72 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.02 2.72 10.72 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.58 1.12 3.22 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.86 2.72 2.40 3.22 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.56 3.04 14.50 3.04 14.50 4.54 14.18 4.54 14.18 3.77
                 13.11 3.77 13.11 4.54 12.78 4.54 12.78 3.45 14.18 3.45
                 14.18 2.24 12.78 2.24 12.78 1.22 13.10 1.22 13.10 1.92
                 14.18 1.92 14.18 1.22 14.50 1.22 14.50 2.72 14.56 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  14.72 0.90 13.80 0.90 13.80 1.54 13.48 1.54 13.48 0.90
                 8.88 0.90 8.88 1.54 8.56 1.54 8.56 0.90 2.58 0.90 2.58 1.54
                 2.26 1.54 2.26 0.90 0.00 0.90 0.00 -0.90 14.72 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  14.72 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.62 1.32 4.62
                 1.32 4.86 7.30 4.86 7.30 4.62 7.62 4.62 7.62 4.86 13.48 4.86
                 13.48 4.21 13.80 4.21 13.80 4.86 14.72 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  13.79 2.98 12.42 2.98 12.42 4.54 8.68 4.54 8.68 2.94 9.00 2.94
                 9.00 4.22 12.10 4.22 12.10 1.22 12.42 1.22 12.42 2.66
                 13.79 2.66 ;
        POLYGON  11.78 2.50 11.46 2.50 11.46 2.18 8.32 2.18 8.32 4.30 6.60 4.30
                 6.60 3.98 8.00 3.98 8.00 2.18 6.48 2.18 6.48 1.22 6.80 1.22
                 6.80 1.86 11.78 1.86 ;
        RECT  9.24 1.22 11.72 1.54 ;
        POLYGON  10.92 3.90 9.38 3.90 9.38 2.94 9.70 2.94 9.70 3.58 10.92 3.58 ;
        RECT  7.18 1.22 8.18 1.54 ;
        POLYGON  7.04 3.22 6.12 3.22 6.12 4.54 2.38 4.54 2.38 3.58 2.70 3.58
                 2.70 4.22 5.80 4.22 5.80 1.22 6.12 1.22 6.12 2.90 7.04 2.90 ;
        RECT  2.94 1.22 5.42 1.54 ;
        POLYGON  5.20 2.50 4.88 2.50 4.88 2.18 0.48 2.18 0.48 3.98 2.02 3.98
                 2.02 4.30 0.16 4.30 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 1.86 5.20 1.86 ;
        RECT  3.08 2.94 4.24 3.90 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END exnor3_4

MACRO exnor3_2
    CLASS CORE ;
    FOREIGN exnor3_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.08 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.02 2.72 10.72 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.58 1.12 3.22 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.86 2.72 2.40 3.22 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  13.92 3.04 13.80 3.04 13.80 4.54 13.48 4.54 13.48 1.22
                 13.80 1.22 13.80 2.72 13.92 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  14.08 0.90 13.10 0.90 13.10 1.54 12.78 1.54 12.78 0.90
                 8.88 0.90 8.88 1.54 8.56 1.54 8.56 0.90 2.58 0.90 2.58 1.54
                 2.26 1.54 2.26 0.90 0.00 0.90 0.00 -0.90 14.08 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  14.08 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.62 1.32 4.62
                 1.32 4.86 7.30 4.86 7.30 4.62 7.62 4.62 7.62 4.86 12.78 4.86
                 12.78 3.58 13.10 3.58 13.10 4.86 14.08 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  13.16 2.98 12.42 2.98 12.42 4.54 8.68 4.54 8.68 2.94 9.00 2.94
                 9.00 4.22 12.10 4.22 12.10 1.22 12.42 1.22 12.42 2.66
                 13.16 2.66 ;
        POLYGON  11.78 2.50 11.46 2.50 11.46 2.18 8.32 2.18 8.32 4.30 6.60 4.30
                 6.60 3.98 8.00 3.98 8.00 2.18 6.48 2.18 6.48 1.22 6.80 1.22
                 6.80 1.86 11.78 1.86 ;
        RECT  9.24 1.22 11.72 1.54 ;
        POLYGON  10.92 3.90 9.38 3.90 9.38 2.94 9.70 2.94 9.70 3.58 10.92 3.58 ;
        RECT  7.18 1.22 8.18 1.54 ;
        POLYGON  7.04 3.22 6.12 3.22 6.12 4.54 2.38 4.54 2.38 3.58 2.70 3.58
                 2.70 4.22 5.80 4.22 5.80 1.22 6.12 1.22 6.12 2.90 7.04 2.90 ;
        RECT  2.94 1.22 5.42 1.54 ;
        POLYGON  5.20 2.50 4.88 2.50 4.88 2.18 0.48 2.18 0.48 3.98 2.02 3.98
                 2.02 4.30 0.16 4.30 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 1.86 5.20 1.86 ;
        RECT  3.08 2.94 4.24 3.90 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END exnor3_2

MACRO exnor3_1
    CLASS CORE ;
    FOREIGN exnor3_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.08 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.02 2.72 10.72 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.58 1.12 3.22 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.86 2.72 2.40 3.22 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  13.92 3.04 13.80 3.04 13.80 4.54 13.48 4.54 13.48 1.22
                 13.80 1.22 13.80 2.72 13.92 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  14.08 0.90 13.10 0.90 13.10 1.54 12.78 1.54 12.78 0.90
                 8.88 0.90 8.88 1.54 8.56 1.54 8.56 0.90 2.58 0.90 2.58 1.54
                 2.26 1.54 2.26 0.90 0.00 0.90 0.00 -0.90 14.08 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  14.08 6.66 0.00 6.66 0.00 4.86 1.00 4.86 1.00 4.62 1.32 4.62
                 1.32 4.86 7.30 4.86 7.30 4.62 7.62 4.62 7.62 4.86 12.78 4.86
                 12.78 4.34 13.10 4.34 13.10 4.86 14.08 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  13.16 2.92 12.42 2.92 12.42 4.54 8.68 4.54 8.68 2.94 9.00 2.94
                 9.00 4.22 12.10 4.22 12.10 1.22 12.42 1.22 12.42 2.60
                 13.16 2.60 ;
        POLYGON  11.78 2.50 11.46 2.50 11.46 2.18 8.32 2.18 8.32 4.30 6.60 4.30
                 6.60 3.98 8.00 3.98 8.00 2.18 6.48 2.18 6.48 1.22 6.80 1.22
                 6.80 1.86 11.78 1.86 ;
        RECT  9.24 1.22 11.72 1.54 ;
        POLYGON  10.92 3.90 9.38 3.90 9.38 2.94 9.70 2.94 9.70 3.58 10.92 3.58 ;
        RECT  7.18 1.22 8.18 1.54 ;
        POLYGON  7.04 3.22 6.12 3.22 6.12 4.54 2.38 4.54 2.38 4.22 5.80 4.22
                 5.80 1.22 6.12 1.22 6.12 2.90 7.04 2.90 ;
        RECT  2.94 1.22 5.42 1.54 ;
        POLYGON  5.20 2.50 4.88 2.50 4.88 2.18 0.48 2.18 0.48 3.98 2.02 3.98
                 2.02 4.30 0.16 4.30 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 1.86 5.20 1.86 ;
        RECT  3.08 2.94 4.24 3.90 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END exnor3_1

MACRO exnor2_4
    CLASS CORE ;
    FOREIGN exnor2_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.32 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.96 2.30 2.40 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.32  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.34 1.12 3.04 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.16 3.04 8.12 3.04 8.12 4.54 7.80 4.54 7.80 3.88 6.72 3.88
                 6.72 4.54 6.40 4.54 6.40 3.56 7.80 3.56 7.80 2.16 6.40 2.16
                 6.40 1.22 6.72 1.22 6.72 1.84 7.80 1.84 7.80 1.22 8.12 1.22
                 8.12 2.72 8.16 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 0.90 7.42 0.90 7.42 1.46 7.10 1.46 7.10 0.90 1.32 0.90
                 1.32 1.14 1.00 1.14 1.00 0.90 0.00 0.90 0.00 -0.90 8.32 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.22 2.58 4.22
                 2.58 4.86 7.10 4.86 7.10 4.21 7.42 4.21 7.42 4.86 8.32 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  6.78 2.98 6.04 2.98 6.04 4.54 5.72 4.54 5.72 1.54 2.38 1.54
                 2.38 1.22 6.04 1.22 6.04 2.66 6.78 2.66 ;
        RECT  2.94 4.22 5.34 4.54 ;
        POLYGON  5.12 3.90 0.50 3.90 0.50 4.54 0.18 4.54 0.18 3.90 0.16 3.90
                 0.16 1.46 2.02 1.46 2.02 1.78 0.48 1.78 0.48 3.58 4.80 3.58
                 4.80 2.34 5.12 2.34 ;
        RECT  3.08 1.86 4.08 2.18 ;
        RECT  0.88 4.22 1.88 4.54 ;
    END
END exnor2_4

MACRO exnor2_2
    CLASS CORE ;
    FOREIGN exnor2_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.96 2.30 2.40 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.32  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.34 1.12 3.04 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.52 3.04 7.42 3.04 7.42 4.54 7.10 4.54 7.10 1.64 7.42 1.64
                 7.42 2.72 7.52 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 0.90 6.72 0.90 6.72 1.44 6.40 1.44 6.40 0.90 1.32 0.90
                 1.32 1.14 1.00 1.14 1.00 0.90 0.00 0.90 0.00 -0.90 7.68 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.22 2.58 4.22
                 2.58 4.86 6.40 4.86 6.40 4.22 6.72 4.22 6.72 4.86 7.68 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  6.78 2.99 6.04 2.99 6.04 4.54 5.72 4.54 5.72 1.54 2.38 1.54
                 2.38 1.22 6.04 1.22 6.04 2.67 6.78 2.67 ;
        RECT  2.94 4.22 5.34 4.54 ;
        POLYGON  5.12 3.90 0.50 3.90 0.50 4.54 0.18 4.54 0.18 3.90 0.16 3.90
                 0.16 1.46 2.02 1.46 2.02 1.78 0.48 1.78 0.48 3.58 4.80 3.58
                 4.80 2.34 5.12 2.34 ;
        RECT  3.08 1.86 4.08 2.18 ;
        RECT  0.88 4.22 1.88 4.54 ;
    END
END exnor2_2

MACRO exnor2_1
    CLASS CORE ;
    FOREIGN exnor2_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.96 2.30 2.40 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.32  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.34 1.12 3.04 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.52 3.04 7.42 3.04 7.42 4.30 7.10 4.30 7.10 1.22 7.42 1.22
                 7.42 2.72 7.52 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 0.90 6.72 0.90 6.72 1.54 6.40 1.54 6.40 0.90 1.32 0.90
                 1.32 1.14 1.00 1.14 1.00 0.90 0.00 0.90 0.00 -0.90 7.68 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 6.66 0.00 6.66 0.00 4.86 2.26 4.86 2.26 4.22 2.58 4.22
                 2.58 4.86 6.40 4.86 6.40 3.98 6.72 3.98 6.72 4.86 7.68 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  6.78 3.16 6.04 3.16 6.04 4.54 5.72 4.54 5.72 1.54 2.38 1.54
                 2.38 1.22 6.04 1.22 6.04 2.84 6.78 2.84 ;
        RECT  2.94 4.22 5.34 4.54 ;
        POLYGON  5.12 3.90 0.50 3.90 0.50 4.54 0.18 4.54 0.18 3.90 0.16 3.90
                 0.16 1.46 2.02 1.46 2.02 1.78 0.48 1.78 0.48 3.58 4.80 3.58
                 4.80 2.34 5.12 2.34 ;
        RECT  3.08 1.86 4.08 2.18 ;
        RECT  0.88 4.22 1.88 4.54 ;
    END
END exnor2_1

MACRO dffpsqb_4
    CLASS CORE ;
    FOREIGN dffpsqb_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.20 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.51  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.25 2.92 9.44 2.92 9.44 3.04 9.12 3.04 9.12 2.60 10.25 2.60 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.44 2.93 3.04 2.93 3.04 3.04 2.72 3.04 2.72 2.61 3.44 2.61 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  18.93 4.54 18.61 4.54 18.61 3.04 17.53 3.04 17.53 4.54
                 17.21 4.54 17.21 1.22 17.53 1.22 17.53 2.72 18.61 2.72
                 18.61 1.22 18.93 1.22 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.99  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.76 3.46 1.14 3.46 1.14 3.14 1.44 3.14 1.44 2.72 1.76 2.72 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  19.20 0.90 18.23 0.90 18.23 1.54 17.91 1.54 17.91 0.90
                 14.73 0.90 14.73 1.54 14.41 1.54 14.41 0.90 7.12 0.90
                 7.12 1.48 6.80 1.48 6.80 0.90 2.86 0.90 2.86 1.28 2.54 1.28
                 2.54 0.90 0.00 0.90 0.00 -0.90 19.20 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  19.20 6.66 0.00 6.66 0.00 4.86 2.54 4.86 2.54 4.60 2.86 4.60
                 2.86 4.86 7.36 4.86 7.36 3.74 7.68 3.74 7.68 4.86 9.75 4.86
                 9.75 4.36 10.07 4.36 10.07 4.86 13.37 4.86 13.37 4.60
                 13.69 4.60 13.69 4.86 15.51 4.86 15.51 3.96 15.83 3.96
                 15.83 4.86 17.91 4.86 17.91 3.58 18.23 3.58 18.23 4.86
                 19.20 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  16.89 3.18 16.71 3.18 16.71 4.54 16.39 4.54 16.39 3.18
                 15.49 3.18 15.49 3.64 14.07 3.64 14.07 3.32 15.17 3.32
                 15.17 2.86 16.57 2.86 16.57 1.54 16.49 1.54 16.49 1.22
                 16.89 1.22 ;
        POLYGON  16.17 2.47 15.85 2.47 15.85 2.28 12.23 2.28 12.23 4.54
                 11.91 4.54 11.91 2.02 11.77 1.88 11.77 1.22 12.09 1.22
                 12.09 1.74 12.31 1.96 16.17 1.96 ;
        RECT  15.11 1.22 16.11 1.54 ;
        RECT  12.69 3.96 15.07 4.28 ;
        RECT  12.47 1.22 14.03 1.54 ;
        POLYGON  11.53 4.04 9.89 4.04 9.89 3.68 9.37 3.68 9.37 4.32 9.05 4.32
                 9.05 3.36 10.21 3.36 10.21 3.72 11.53 3.72 ;
        RECT  8.72 1.22 11.39 1.54 ;
        POLYGON  10.93 3.40 10.53 3.40 10.53 3.08 10.61 3.08 10.61 2.18
                 8.08 2.18 8.08 1.86 10.93 1.86 ;
        POLYGON  8.51 4.48 8.19 4.48 8.19 2.82 5.36 2.82 5.36 2.26 5.68 2.26
                 5.68 2.50 7.44 2.50 7.44 1.22 8.38 1.22 8.38 1.54 7.76 1.54
                 7.76 2.50 8.51 2.50 ;
        RECT  5.83 3.46 6.87 3.78 ;
        POLYGON  6.51 4.54 3.18 4.54 3.18 4.28 2.16 4.28 2.16 4.54 0.46 4.54
                 0.46 1.22 0.78 1.22 0.78 4.22 1.84 4.22 1.84 3.96 3.50 3.96
                 3.50 4.22 6.51 4.22 ;
        RECT  5.42 1.22 6.42 1.54 ;
        POLYGON  5.45 3.90 4.72 3.90 4.72 2.18 2.49 2.18 2.49 2.38 2.17 2.38
                 2.17 1.86 4.72 1.86 4.72 1.22 5.04 1.22 5.04 3.58 5.45 3.58 ;
        RECT  3.24 1.22 4.34 1.54 ;
        RECT  3.24 3.32 4.34 3.64 ;
        RECT  1.16 1.22 2.16 1.54 ;
    END
END dffpsqb_4

MACRO dffpsqb_2
    CLASS CORE ;
    FOREIGN dffpsqb_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.56 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.51  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.25 2.92 9.44 2.92 9.44 3.04 9.12 3.04 9.12 2.60 10.25 2.60 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.44 2.93 3.04 2.93 3.04 3.04 2.72 3.04 2.72 2.61 3.44 2.61 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  18.40 3.04 18.19 3.04 18.19 4.54 17.87 4.54 17.87 1.39
                 18.19 1.39 18.19 2.72 18.40 2.72 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.99  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.76 3.46 1.14 3.46 1.14 3.14 1.44 3.14 1.44 2.72 1.76 2.72 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  18.56 0.90 17.49 0.90 17.49 1.49 17.17 1.49 17.17 0.90
                 14.73 0.90 14.73 1.54 14.41 1.54 14.41 0.90 7.12 0.90
                 7.12 1.48 6.80 1.48 6.80 0.90 0.00 0.90 0.00 -0.90 18.56 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  18.56 6.66 0.00 6.66 0.00 4.86 2.54 4.86 2.54 4.60 2.86 4.60
                 2.86 4.86 7.36 4.86 7.36 3.74 7.68 3.74 7.68 4.86 9.75 4.86
                 9.75 4.36 10.07 4.36 10.07 4.86 13.37 4.86 13.37 4.60
                 13.69 4.60 13.69 4.86 15.51 4.86 15.51 3.96 15.83 3.96
                 15.83 4.86 17.17 4.86 17.17 3.59 17.49 3.59 17.49 4.86
                 18.56 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  17.00 2.46 16.81 2.46 16.81 3.18 16.71 3.18 16.71 4.54
                 16.39 4.54 16.39 3.18 15.49 3.18 15.49 3.64 14.07 3.64
                 14.07 3.32 15.17 3.32 15.17 2.86 16.49 2.86 16.49 1.22
                 16.81 1.22 16.81 2.13 17.00 2.13 ;
        POLYGON  16.17 2.47 15.85 2.47 15.85 2.28 12.23 2.28 12.23 4.54
                 11.91 4.54 11.91 2.02 11.77 1.88 11.77 1.22 12.09 1.22
                 12.09 1.74 12.31 1.96 16.17 1.96 ;
        RECT  15.11 1.22 16.11 1.54 ;
        RECT  12.69 3.96 15.07 4.28 ;
        RECT  12.47 1.22 14.03 1.54 ;
        POLYGON  11.53 4.04 9.89 4.04 9.89 3.68 9.37 3.68 9.37 4.32 9.05 4.32
                 9.05 3.36 10.21 3.36 10.21 3.72 11.53 3.72 ;
        RECT  8.72 1.22 11.39 1.54 ;
        POLYGON  10.93 3.40 10.53 3.40 10.53 3.08 10.61 3.08 10.61 2.18
                 8.08 2.18 8.08 1.86 10.93 1.86 ;
        POLYGON  8.51 4.48 8.19 4.48 8.19 2.82 5.36 2.82 5.36 2.26 5.68 2.26
                 5.68 2.50 7.44 2.50 7.44 1.22 8.38 1.22 8.38 1.54 7.76 1.54
                 7.76 2.50 8.51 2.50 ;
        RECT  5.83 3.46 6.87 3.78 ;
        POLYGON  6.51 4.54 3.18 4.54 3.18 4.28 2.16 4.28 2.16 4.54 0.46 4.54
                 0.46 1.22 0.78 1.22 0.78 4.22 1.84 4.22 1.84 3.96 3.50 3.96
                 3.50 4.22 6.51 4.22 ;
        RECT  5.42 1.22 6.42 1.54 ;
        POLYGON  5.45 3.90 4.72 3.90 4.72 2.18 2.49 2.18 2.49 2.38 2.17 2.38
                 2.17 1.86 4.72 1.86 4.72 1.22 5.04 1.22 5.04 3.58 5.45 3.58 ;
        RECT  3.24 1.22 4.34 1.54 ;
        RECT  3.24 3.32 4.34 3.64 ;
        RECT  1.16 1.22 2.16 1.54 ;
    END
END dffpsqb_2

MACRO dffpsqb_1
    CLASS CORE ;
    FOREIGN dffpsqb_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.56 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.51  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.25 2.92 9.44 2.92 9.44 3.04 9.12 3.04 9.12 2.60 10.25 2.60 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.44 2.93 3.04 2.93 3.04 3.04 2.72 3.04 2.72 2.61 3.44 2.61 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  18.40 3.04 18.19 3.04 18.19 4.30 17.87 4.30 17.87 1.22
                 18.19 1.22 18.19 2.72 18.40 2.72 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.99  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.76 3.46 1.14 3.46 1.14 3.14 1.44 3.14 1.44 2.72 1.76 2.72 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  18.56 0.90 17.49 0.90 17.49 1.55 17.17 1.55 17.17 0.90
                 14.73 0.90 14.73 1.54 14.41 1.54 14.41 0.90 7.12 0.90
                 7.12 1.48 6.80 1.48 6.80 0.90 2.86 0.90 2.86 1.28 2.54 1.28
                 2.54 0.90 0.00 0.90 0.00 -0.90 18.56 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  18.56 6.66 0.00 6.66 0.00 4.86 2.54 4.86 2.54 4.60 2.86 4.60
                 2.86 4.86 7.36 4.86 7.36 3.74 7.68 3.74 7.68 4.86 9.75 4.86
                 9.75 4.36 10.07 4.36 10.07 4.86 13.37 4.86 13.37 4.60
                 13.69 4.60 13.69 4.86 15.51 4.86 15.51 3.96 15.83 3.96
                 15.83 4.86 17.17 4.86 17.17 3.98 17.49 3.98 17.49 4.86
                 18.56 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  16.99 2.46 16.81 2.46 16.81 3.18 16.71 3.18 16.71 4.54
                 16.39 4.54 16.39 3.18 15.49 3.18 15.49 3.64 14.07 3.64
                 14.07 3.32 15.17 3.32 15.17 2.86 16.49 2.86 16.49 1.22
                 16.81 1.22 16.81 2.14 16.99 2.14 ;
        POLYGON  16.17 2.47 15.85 2.47 15.85 2.28 12.23 2.28 12.23 4.54
                 11.91 4.54 11.91 2.02 11.77 1.88 11.77 1.22 12.09 1.22
                 12.09 1.74 12.31 1.96 16.17 1.96 ;
        RECT  15.11 1.22 16.11 1.54 ;
        RECT  12.69 3.96 15.07 4.28 ;
        RECT  12.47 1.22 14.03 1.54 ;
        POLYGON  11.53 4.04 9.89 4.04 9.89 3.68 9.37 3.68 9.37 4.32 9.05 4.32
                 9.05 3.36 10.21 3.36 10.21 3.72 11.53 3.72 ;
        RECT  8.72 1.22 11.39 1.54 ;
        POLYGON  10.93 3.40 10.53 3.40 10.53 3.08 10.61 3.08 10.61 2.18
                 8.08 2.18 8.08 1.86 10.93 1.86 ;
        POLYGON  8.51 4.48 8.19 4.48 8.19 2.82 5.36 2.82 5.36 2.26 5.68 2.26
                 5.68 2.50 7.44 2.50 7.44 1.22 8.38 1.22 8.38 1.54 7.76 1.54
                 7.76 2.50 8.51 2.50 ;
        RECT  5.83 3.46 6.87 3.78 ;
        POLYGON  6.51 4.54 3.18 4.54 3.18 4.28 2.16 4.28 2.16 4.54 0.46 4.54
                 0.46 1.22 0.78 1.22 0.78 4.22 1.84 4.22 1.84 3.96 3.50 3.96
                 3.50 4.22 6.51 4.22 ;
        RECT  5.42 1.22 6.42 1.54 ;
        POLYGON  5.45 3.90 4.72 3.90 4.72 2.18 2.49 2.18 2.49 2.38 2.17 2.38
                 2.17 1.86 4.72 1.86 4.72 1.22 5.04 1.22 5.04 3.58 5.45 3.58 ;
        RECT  3.24 1.22 4.34 1.54 ;
        RECT  3.24 3.32 4.34 3.64 ;
        RECT  1.16 1.22 2.16 1.54 ;
    END
END dffpsqb_1

MACRO dffpsq_4
    CLASS CORE ;
    FOREIGN dffpsq_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.20 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.51  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.25 2.92 9.44 2.92 9.44 3.04 9.12 3.04 9.12 2.60 10.25 2.60 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.44 2.93 3.04 2.93 3.04 3.04 2.72 3.04 2.72 2.61 3.44 2.61 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  18.89 4.54 18.57 4.54 18.57 3.04 17.49 3.04 17.49 4.54
                 17.17 4.54 17.17 1.22 17.49 1.22 17.49 2.72 18.57 2.72
                 18.57 1.22 18.89 1.22 ;
        END
    END q
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.99  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.76 3.46 1.14 3.46 1.14 3.14 1.44 3.14 1.44 2.72 1.76 2.72 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  19.20 0.90 18.19 0.90 18.19 1.54 17.87 1.54 17.87 0.90
                 14.73 0.90 14.73 1.54 14.41 1.54 14.41 0.90 7.12 0.90
                 7.12 1.48 6.80 1.48 6.80 0.90 2.86 0.90 2.86 1.28 2.54 1.28
                 2.54 0.90 0.00 0.90 0.00 -0.90 19.20 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  19.20 6.66 0.00 6.66 0.00 4.86 2.54 4.86 2.54 4.60 2.86 4.60
                 2.86 4.86 7.36 4.86 7.36 3.74 7.68 3.74 7.68 4.86 9.75 4.86
                 9.75 4.36 10.07 4.36 10.07 4.86 13.37 4.86 13.37 4.60
                 13.69 4.60 13.69 4.86 15.51 4.86 15.51 3.96 15.83 3.96
                 15.83 4.86 17.87 4.86 17.87 3.58 18.19 3.58 18.19 4.86
                 19.20 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  16.81 3.18 16.71 3.18 16.71 4.54 16.39 4.54 16.39 3.18
                 15.49 3.18 15.49 3.64 14.07 3.64 14.07 3.32 15.17 3.32
                 15.17 2.86 16.49 2.86 16.49 1.22 16.81 1.22 ;
        POLYGON  16.17 2.47 15.85 2.47 15.85 2.28 12.23 2.28 12.23 4.54
                 11.91 4.54 11.91 2.02 11.77 1.88 11.77 1.22 12.09 1.22
                 12.09 1.74 12.31 1.96 16.17 1.96 ;
        RECT  15.11 1.22 16.11 1.54 ;
        RECT  12.69 3.96 15.07 4.28 ;
        RECT  12.47 1.22 14.03 1.54 ;
        POLYGON  11.53 4.04 9.89 4.04 9.89 3.68 9.37 3.68 9.37 4.32 9.05 4.32
                 9.05 3.36 10.21 3.36 10.21 3.72 11.53 3.72 ;
        RECT  8.72 1.22 11.39 1.54 ;
        POLYGON  10.93 3.40 10.53 3.40 10.53 3.08 10.61 3.08 10.61 2.18
                 8.08 2.18 8.08 1.86 10.93 1.86 ;
        POLYGON  8.51 4.48 8.19 4.48 8.19 2.82 5.36 2.82 5.36 2.26 5.68 2.26
                 5.68 2.50 7.44 2.50 7.44 1.22 8.38 1.22 8.38 1.54 7.76 1.54
                 7.76 2.50 8.51 2.50 ;
        RECT  5.83 3.46 6.87 3.78 ;
        POLYGON  6.51 4.54 3.18 4.54 3.18 4.28 2.16 4.28 2.16 4.54 0.46 4.54
                 0.46 1.22 0.78 1.22 0.78 4.22 1.84 4.22 1.84 3.96 3.50 3.96
                 3.50 4.22 6.51 4.22 ;
        RECT  5.42 1.22 6.42 1.54 ;
        POLYGON  5.45 3.90 4.72 3.90 4.72 2.18 2.49 2.18 2.49 2.38 2.17 2.38
                 2.17 1.86 4.72 1.86 4.72 1.22 5.04 1.22 5.04 3.58 5.45 3.58 ;
        RECT  3.24 1.22 4.34 1.54 ;
        RECT  3.24 3.32 4.34 3.64 ;
        RECT  1.16 1.22 2.16 1.54 ;
    END
END dffpsq_4

MACRO dffpsq_2
    CLASS CORE ;
    FOREIGN dffpsq_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.56 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.51  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.25 2.92 9.44 2.92 9.44 3.04 9.12 3.04 9.12 2.60 10.25 2.60 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.44 2.93 3.04 2.93 3.04 3.04 2.72 3.04 2.72 2.61 3.44 2.61 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  18.40 3.04 18.19 3.04 18.19 4.54 17.87 4.54 17.87 1.39
                 18.19 1.39 18.19 2.72 18.40 2.72 ;
        END
    END q
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.99  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.76 3.46 1.14 3.46 1.14 3.14 1.44 3.14 1.44 2.72 1.76 2.72 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  18.56 0.90 17.49 0.90 17.49 1.49 17.17 1.49 17.17 0.90
                 14.73 0.90 14.73 1.54 14.41 1.54 14.41 0.90 7.12 0.90
                 7.12 1.48 6.80 1.48 6.80 0.90 0.00 0.90 0.00 -0.90 18.56 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  18.56 6.66 0.00 6.66 0.00 4.86 2.54 4.86 2.54 4.60 2.86 4.60
                 2.86 4.86 7.36 4.86 7.36 3.74 7.68 3.74 7.68 4.86 9.75 4.86
                 9.75 4.36 10.07 4.36 10.07 4.86 13.37 4.86 13.37 4.60
                 13.69 4.60 13.69 4.86 15.51 4.86 15.51 3.96 15.83 3.96
                 15.83 4.86 17.17 4.86 17.17 3.59 17.49 3.59 17.49 4.86
                 18.56 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  16.81 3.18 16.71 3.18 16.71 4.54 16.39 4.54 16.39 3.18
                 15.49 3.18 15.49 3.64 14.07 3.64 14.07 3.32 15.17 3.32
                 15.17 2.86 16.49 2.86 16.49 1.22 16.81 1.22 ;
        POLYGON  16.17 2.47 15.85 2.47 15.85 2.28 12.23 2.28 12.23 4.54
                 11.91 4.54 11.91 2.02 11.77 1.88 11.77 1.22 12.09 1.22
                 12.09 1.74 12.31 1.96 16.17 1.96 ;
        RECT  15.11 1.22 16.11 1.54 ;
        RECT  12.69 3.96 15.07 4.28 ;
        RECT  12.47 1.22 14.03 1.54 ;
        POLYGON  11.53 4.04 9.89 4.04 9.89 3.68 9.37 3.68 9.37 4.32 9.05 4.32
                 9.05 3.36 10.21 3.36 10.21 3.72 11.53 3.72 ;
        RECT  8.72 1.22 11.39 1.54 ;
        POLYGON  10.93 3.40 10.53 3.40 10.53 3.08 10.61 3.08 10.61 2.18
                 8.08 2.18 8.08 1.86 10.93 1.86 ;
        POLYGON  8.51 4.48 8.19 4.48 8.19 2.82 5.36 2.82 5.36 2.26 5.68 2.26
                 5.68 2.50 7.44 2.50 7.44 1.22 8.38 1.22 8.38 1.54 7.76 1.54
                 7.76 2.50 8.51 2.50 ;
        RECT  5.83 3.46 6.87 3.78 ;
        POLYGON  6.51 4.54 3.18 4.54 3.18 4.28 2.16 4.28 2.16 4.54 0.46 4.54
                 0.46 1.22 0.78 1.22 0.78 4.22 1.84 4.22 1.84 3.96 3.50 3.96
                 3.50 4.22 6.51 4.22 ;
        RECT  5.42 1.22 6.42 1.54 ;
        POLYGON  5.45 3.90 4.72 3.90 4.72 2.18 2.49 2.18 2.49 2.38 2.17 2.38
                 2.17 1.86 4.72 1.86 4.72 1.22 5.04 1.22 5.04 3.58 5.45 3.58 ;
        RECT  3.24 1.22 4.34 1.54 ;
        RECT  3.24 3.32 4.34 3.64 ;
        RECT  1.16 1.22 2.16 1.54 ;
    END
END dffpsq_2

MACRO dffpsq_1
    CLASS CORE ;
    FOREIGN dffpsq_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.56 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.51  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.25 2.92 9.44 2.92 9.44 3.04 9.12 3.04 9.12 2.60 10.25 2.60 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.44 2.93 3.04 2.93 3.04 3.04 2.72 3.04 2.72 2.61 3.44 2.61 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  18.40 3.04 18.19 3.04 18.19 4.30 17.87 4.30 17.87 1.22
                 18.19 1.22 18.19 2.72 18.40 2.72 ;
        END
    END q
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.99  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.76 3.46 1.14 3.46 1.14 3.14 1.44 3.14 1.44 2.72 1.76 2.72 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  18.56 0.90 17.49 0.90 17.49 1.55 17.17 1.55 17.17 0.90
                 14.73 0.90 14.73 1.54 14.41 1.54 14.41 0.90 7.12 0.90
                 7.12 1.48 6.80 1.48 6.80 0.90 2.86 0.90 2.86 1.28 2.54 1.28
                 2.54 0.90 0.00 0.90 0.00 -0.90 18.56 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  18.56 6.66 0.00 6.66 0.00 4.86 2.54 4.86 2.54 4.60 2.86 4.60
                 2.86 4.86 7.36 4.86 7.36 3.74 7.68 3.74 7.68 4.86 9.75 4.86
                 9.75 4.36 10.07 4.36 10.07 4.86 13.37 4.86 13.37 4.60
                 13.69 4.60 13.69 4.86 15.51 4.86 15.51 3.96 15.83 3.96
                 15.83 4.86 17.17 4.86 17.17 3.98 17.49 3.98 17.49 4.86
                 18.56 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  16.81 3.18 16.71 3.18 16.71 4.54 16.39 4.54 16.39 3.18
                 15.49 3.18 15.49 3.64 14.07 3.64 14.07 3.32 15.17 3.32
                 15.17 2.86 16.49 2.86 16.49 1.22 16.81 1.22 ;
        POLYGON  16.17 2.47 15.85 2.47 15.85 2.28 12.23 2.28 12.23 4.54
                 11.91 4.54 11.91 2.02 11.77 1.88 11.77 1.22 12.09 1.22
                 12.09 1.74 12.31 1.96 16.17 1.96 ;
        RECT  15.11 1.22 16.11 1.54 ;
        RECT  12.69 3.96 15.07 4.28 ;
        RECT  12.47 1.22 14.03 1.54 ;
        POLYGON  11.53 4.04 9.89 4.04 9.89 3.68 9.37 3.68 9.37 4.32 9.05 4.32
                 9.05 3.36 10.21 3.36 10.21 3.72 11.53 3.72 ;
        RECT  8.72 1.22 11.39 1.54 ;
        POLYGON  10.93 3.40 10.53 3.40 10.53 3.08 10.61 3.08 10.61 2.18
                 8.08 2.18 8.08 1.86 10.93 1.86 ;
        POLYGON  8.51 4.48 8.19 4.48 8.19 2.82 5.36 2.82 5.36 2.26 5.68 2.26
                 5.68 2.50 7.44 2.50 7.44 1.22 8.38 1.22 8.38 1.54 7.76 1.54
                 7.76 2.50 8.51 2.50 ;
        RECT  5.83 3.46 6.87 3.78 ;
        POLYGON  6.51 4.54 3.18 4.54 3.18 4.28 2.16 4.28 2.16 4.54 0.46 4.54
                 0.46 1.22 0.78 1.22 0.78 4.22 1.84 4.22 1.84 3.96 3.50 3.96
                 3.50 4.22 6.51 4.22 ;
        RECT  5.42 1.22 6.42 1.54 ;
        POLYGON  5.45 3.90 4.72 3.90 4.72 2.18 2.49 2.18 2.49 2.38 2.17 2.38
                 2.17 1.86 4.72 1.86 4.72 1.22 5.04 1.22 5.04 3.58 5.45 3.58 ;
        RECT  3.24 1.22 4.34 1.54 ;
        RECT  3.24 3.32 4.34 3.64 ;
        RECT  1.16 1.22 2.16 1.54 ;
    END
END dffpsq_1

MACRO dffps_4
    CLASS CORE ;
    FOREIGN dffps_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.76 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.51  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.25 2.92 9.44 2.92 9.44 3.04 9.12 3.04 9.12 2.60 10.25 2.60 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.44 2.93 3.04 2.93 3.04 3.04 2.72 3.04 2.72 2.61 3.44 2.61 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  19.38 3.25 17.65 3.25 17.65 2.93 18.72 2.93 18.72 2.71
                 19.06 2.71 19.06 1.54 17.17 1.54 17.17 1.22 19.38 1.22 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  21.60 3.04 21.48 3.04 21.48 4.53 19.74 4.53 19.74 4.21
                 21.16 4.21 21.16 1.90 19.74 1.90 19.74 1.58 21.48 1.58
                 21.48 2.72 21.60 2.72 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.99  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.76 3.46 1.14 3.46 1.14 3.14 1.44 3.14 1.44 2.72 1.76 2.72 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.76 0.90 14.73 0.90 14.73 1.54 14.41 1.54 14.41 0.90
                 7.12 0.90 7.12 1.48 6.80 1.48 6.80 0.90 2.86 0.90 2.86 1.28
                 2.54 1.28 2.54 0.90 0.00 0.90 0.00 -0.90 21.76 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.76 6.66 0.00 6.66 0.00 4.86 2.54 4.86 2.54 4.60 2.86 4.60
                 2.86 4.86 7.36 4.86 7.36 3.74 7.68 3.74 7.68 4.86 9.75 4.86
                 9.75 4.36 10.07 4.36 10.07 4.86 13.37 4.86 13.37 4.60
                 13.69 4.60 13.69 4.86 15.51 4.86 15.51 3.96 15.83 3.96
                 15.83 4.86 18.29 4.86 18.29 4.79 18.71 4.79 18.71 4.86
                 21.76 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.76 3.89 18.13 3.89 18.13 4.32 16.39 4.32 16.39 3.18
                 15.49 3.18 15.49 3.64 14.07 3.64 14.07 3.32 15.17 3.32
                 15.17 2.86 16.49 2.86 16.49 1.22 16.81 1.22 16.81 3.18
                 16.71 3.18 16.71 4.00 17.81 4.00 17.81 3.57 20.44 3.57
                 20.44 2.33 20.76 2.33 ;
        POLYGON  16.17 2.47 15.85 2.47 15.85 2.28 12.23 2.28 12.23 4.54
                 11.91 4.54 11.91 2.02 11.77 1.88 11.77 1.22 12.09 1.22
                 12.09 1.74 12.31 1.96 16.17 1.96 ;
        RECT  15.11 1.22 16.11 1.54 ;
        RECT  12.69 3.96 15.07 4.28 ;
        RECT  12.47 1.22 14.03 1.54 ;
        POLYGON  11.53 4.04 9.89 4.04 9.89 3.68 9.05 3.68 9.05 3.36 10.21 3.36
                 10.21 3.72 11.53 3.72 ;
        RECT  8.72 1.22 11.39 1.54 ;
        POLYGON  10.93 3.40 10.53 3.40 10.53 3.08 10.61 3.08 10.61 2.18
                 8.08 2.18 8.08 1.86 10.93 1.86 ;
        POLYGON  8.51 3.90 8.19 3.90 8.19 2.82 5.36 2.82 5.36 2.26 5.68 2.26
                 5.68 2.50 7.44 2.50 7.44 1.22 8.38 1.22 8.38 1.54 7.76 1.54
                 7.76 2.50 8.51 2.50 ;
        RECT  5.83 3.46 6.87 3.78 ;
        POLYGON  6.51 4.54 3.18 4.54 3.18 4.28 2.16 4.28 2.16 4.54 0.46 4.54
                 0.46 1.22 0.78 1.22 0.78 4.22 1.84 4.22 1.84 3.96 3.50 3.96
                 3.50 4.22 6.51 4.22 ;
        RECT  5.42 1.22 6.42 1.54 ;
        POLYGON  5.45 3.90 4.72 3.90 4.72 2.18 2.49 2.18 2.49 2.38 2.17 2.38
                 2.17 1.86 4.72 1.86 4.72 1.22 5.04 1.22 5.04 3.58 5.45 3.58 ;
        RECT  3.24 1.22 4.34 1.54 ;
        RECT  3.24 3.32 4.34 3.64 ;
        RECT  1.16 1.22 2.16 1.54 ;
    END
END dffps_4

MACRO dffps_2
    CLASS CORE ;
    FOREIGN dffps_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.20 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.51  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.25 2.92 9.44 2.92 9.44 3.04 9.12 3.04 9.12 2.60 10.25 2.60 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.44 2.93 3.04 2.93 3.04 3.04 2.72 3.04 2.72 2.61 3.44 2.61 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  17.76 3.04 17.49 3.04 17.49 3.42 17.17 3.42 17.17 1.22
                 17.49 1.22 17.49 2.72 17.76 2.72 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  19.04 4.32 18.57 4.32 18.57 4.00 18.72 4.00 18.72 1.55
                 18.57 1.55 18.57 1.23 19.04 1.23 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.99  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.76 3.46 1.14 3.46 1.14 3.14 1.44 3.14 1.44 2.72 1.76 2.72 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  19.20 0.90 18.19 0.90 18.19 1.35 17.87 1.35 17.87 0.90
                 14.73 0.90 14.73 1.54 14.41 1.54 14.41 0.90 7.12 0.90
                 7.12 1.48 6.80 1.48 6.80 0.90 2.86 0.90 2.86 1.28 2.54 1.28
                 2.54 0.90 0.00 0.90 0.00 -0.90 19.20 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  19.20 6.66 0.00 6.66 0.00 4.86 2.54 4.86 2.54 4.60 2.86 4.60
                 2.86 4.86 7.36 4.86 7.36 3.74 7.68 3.74 7.68 4.86 9.75 4.86
                 9.75 4.36 10.07 4.36 10.07 4.86 13.37 4.86 13.37 4.60
                 13.69 4.60 13.69 4.86 15.51 4.86 15.51 3.96 15.83 3.96
                 15.83 4.86 19.20 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  18.40 3.68 18.13 3.68 18.13 4.54 16.39 4.54 16.39 3.18
                 15.49 3.18 15.49 3.64 14.07 3.64 14.07 3.32 15.17 3.32
                 15.17 2.86 16.49 2.86 16.49 1.22 16.81 1.22 16.81 3.18
                 16.71 3.18 16.71 4.22 17.81 4.22 17.81 3.36 18.08 3.36
                 18.08 2.46 18.03 2.46 18.03 2.14 18.40 2.14 ;
        POLYGON  16.17 2.47 15.85 2.47 15.85 2.28 12.23 2.28 12.23 4.54
                 11.91 4.54 11.91 2.02 11.77 1.88 11.77 1.22 12.09 1.22
                 12.09 1.74 12.31 1.96 16.17 1.96 ;
        RECT  15.11 1.22 16.11 1.54 ;
        RECT  12.69 3.96 15.07 4.28 ;
        RECT  12.47 1.22 14.03 1.54 ;
        POLYGON  11.53 4.04 9.89 4.04 9.89 3.68 9.05 3.68 9.05 3.36 10.21 3.36
                 10.21 3.72 11.53 3.72 ;
        RECT  8.72 1.22 11.39 1.54 ;
        POLYGON  10.93 3.40 10.53 3.40 10.53 3.08 10.61 3.08 10.61 2.18
                 8.08 2.18 8.08 1.86 10.93 1.86 ;
        POLYGON  8.51 3.90 8.19 3.90 8.19 2.82 5.36 2.82 5.36 2.26 5.68 2.26
                 5.68 2.50 7.44 2.50 7.44 1.22 8.38 1.22 8.38 1.54 7.76 1.54
                 7.76 2.50 8.51 2.50 ;
        RECT  5.83 3.46 6.87 3.78 ;
        POLYGON  6.51 4.54 3.18 4.54 3.18 4.28 2.16 4.28 2.16 4.54 0.46 4.54
                 0.46 1.22 0.78 1.22 0.78 4.22 1.84 4.22 1.84 3.96 3.50 3.96
                 3.50 4.22 6.51 4.22 ;
        RECT  5.42 1.22 6.42 1.54 ;
        POLYGON  5.45 3.90 4.72 3.90 4.72 2.18 2.49 2.18 2.49 2.38 2.17 2.38
                 2.17 1.86 4.72 1.86 4.72 1.22 5.04 1.22 5.04 3.58 5.45 3.58 ;
        RECT  3.24 1.22 4.34 1.54 ;
        RECT  3.24 3.32 4.34 3.64 ;
        RECT  1.16 1.22 2.16 1.54 ;
    END
END dffps_2

MACRO dffps_1
    CLASS CORE ;
    FOREIGN dffps_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.20 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.51  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.25 2.92 9.44 2.92 9.44 3.04 9.12 3.04 9.12 2.60 10.25 2.60 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.44 2.93 3.04 2.93 3.04 3.04 2.72 3.04 2.72 2.61 3.44 2.61 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.21  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  17.76 3.04 17.49 3.04 17.49 3.90 17.17 3.90 17.17 1.22
                 17.49 1.22 17.49 2.72 17.76 2.72 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.21  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  19.04 4.32 18.57 4.32 18.57 4.00 18.72 4.00 18.72 1.55
                 18.57 1.55 18.57 1.23 19.04 1.23 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.99  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.76 3.46 1.14 3.46 1.14 3.14 1.44 3.14 1.44 2.72 1.76 2.72 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  19.20 0.90 18.19 0.90 18.19 1.54 17.87 1.54 17.87 0.90
                 14.73 0.90 14.73 1.54 14.41 1.54 14.41 0.90 7.12 0.90
                 7.12 1.48 6.80 1.48 6.80 0.90 2.86 0.90 2.86 1.28 2.54 1.28
                 2.54 0.90 0.00 0.90 0.00 -0.90 19.20 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  19.20 6.66 0.00 6.66 0.00 4.86 2.54 4.86 2.54 4.60 2.86 4.60
                 2.86 4.86 7.36 4.86 7.36 3.74 7.68 3.74 7.68 4.86 9.75 4.86
                 9.75 4.36 10.07 4.36 10.07 4.86 13.37 4.86 13.37 4.60
                 13.69 4.60 13.69 4.86 15.51 4.86 15.51 3.96 15.83 3.96
                 15.83 4.86 19.20 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  18.40 3.68 18.13 3.68 18.13 4.54 16.39 4.54 16.39 3.18
                 15.49 3.18 15.49 3.64 14.07 3.64 14.07 3.32 15.17 3.32
                 15.17 2.86 16.49 2.86 16.49 1.22 16.81 1.22 16.81 3.18
                 16.71 3.18 16.71 4.22 17.81 4.22 17.81 3.36 18.08 3.36
                 18.08 2.46 18.03 2.46 18.03 2.14 18.40 2.14 ;
        POLYGON  16.17 2.47 15.85 2.47 15.85 2.28 12.23 2.28 12.23 4.54
                 11.91 4.54 11.91 2.02 11.77 1.88 11.77 1.22 12.09 1.22
                 12.09 1.74 12.31 1.96 16.17 1.96 ;
        RECT  15.11 1.22 16.11 1.54 ;
        RECT  12.69 3.96 15.07 4.28 ;
        RECT  12.47 1.22 14.03 1.54 ;
        POLYGON  11.53 4.04 9.89 4.04 9.89 3.68 9.05 3.68 9.05 3.36 10.21 3.36
                 10.21 3.72 11.53 3.72 ;
        RECT  8.72 1.22 11.39 1.54 ;
        POLYGON  10.93 3.40 10.53 3.40 10.53 3.08 10.61 3.08 10.61 2.18
                 8.08 2.18 8.08 1.86 10.93 1.86 ;
        POLYGON  8.51 3.90 8.19 3.90 8.19 2.82 5.36 2.82 5.36 2.26 5.68 2.26
                 5.68 2.50 7.44 2.50 7.44 1.22 8.38 1.22 8.38 1.54 7.76 1.54
                 7.76 2.50 8.51 2.50 ;
        RECT  5.83 3.46 6.87 3.78 ;
        POLYGON  6.51 4.54 3.18 4.54 3.18 4.28 2.16 4.28 2.16 4.54 0.46 4.54
                 0.46 1.22 0.78 1.22 0.78 4.22 1.84 4.22 1.84 3.96 3.50 3.96
                 3.50 4.22 6.51 4.22 ;
        RECT  5.42 1.22 6.42 1.54 ;
        POLYGON  5.45 3.90 4.72 3.90 4.72 2.18 2.49 2.18 2.49 2.38 2.17 2.38
                 2.17 1.86 4.72 1.86 4.72 1.22 5.04 1.22 5.04 3.58 5.45 3.58 ;
        RECT  3.24 1.22 4.34 1.54 ;
        RECT  3.24 3.32 4.34 3.64 ;
        RECT  1.16 1.22 2.16 1.54 ;
    END
END dffps_1

MACRO dffprsqb_4
    CLASS CORE ;
    FOREIGN dffprsqb_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.64 2.72 11.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.72 4.64 3.04 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.97  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.96 3.04 20.74 3.04 20.74 4.54 20.42 4.54 20.42 1.22
                 20.74 1.22 20.74 2.72 20.96 2.72 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.12 0.52 3.04 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.28 2.50 3.68 3.06 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  22.40 0.90 21.44 0.90 21.44 1.56 21.12 1.56 21.12 0.90
                 19.86 0.90 19.86 1.54 19.54 1.54 19.54 0.90 16.64 0.90
                 16.64 1.54 16.32 1.54 16.32 0.90 4.20 0.90 4.20 1.54 3.88 1.54
                 3.88 0.90 0.00 0.90 0.00 -0.90 22.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  22.40 6.66 0.00 6.66 0.00 4.86 0.99 4.86 0.99 4.16 1.31 4.16
                 1.31 4.86 5.52 4.86 5.52 4.62 5.84 4.62 5.84 4.86 9.40 4.86
                 9.40 4.16 9.72 4.16 9.72 4.86 11.68 4.86 11.68 4.64 12.00 4.64
                 12.00 4.86 15.32 4.86 15.32 3.94 15.64 3.94 15.64 4.86
                 19.60 4.86 19.60 4.26 19.92 4.26 19.92 4.86 21.12 4.86
                 21.12 3.80 21.44 3.80 21.44 4.86 22.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.10 3.06 18.42 3.06 18.42 3.90 18.10 3.90 18.10 3.06
                 17.02 3.06 17.02 4.54 16.70 4.54 16.70 2.86 15.92 2.86
                 15.92 2.54 17.02 2.54 17.02 2.74 18.78 2.74 18.78 1.22
                 19.10 1.22 19.10 2.74 19.78 2.74 19.78 2.62 20.10 2.62 ;
        POLYGON  19.10 4.54 17.40 4.54 17.40 3.58 17.72 3.58 17.72 4.22
                 19.10 4.22 ;
        POLYGON  18.12 2.42 17.79 2.42 17.79 2.18 14.56 2.18 14.56 2.70
                 14.16 3.10 14.16 4.12 13.84 4.12 13.84 2.96 14.24 2.56
                 14.24 1.22 14.56 1.22 14.56 1.86 18.12 1.86 ;
        RECT  17.02 1.22 18.02 1.54 ;
        POLYGON  16.34 3.62 14.86 3.62 14.86 3.80 14.54 3.80 14.54 3.30
                 16.34 3.30 ;
        RECT  14.94 1.22 15.94 1.54 ;
        RECT  11.30 1.22 13.86 1.54 ;
        POLYGON  13.82 2.44 13.26 2.44 13.26 3.68 12.46 3.68 12.46 3.36
                 12.94 3.36 12.94 2.18 10.66 2.18 10.66 1.54 9.10 1.54
                 9.10 2.38 7.04 2.38 7.04 2.06 8.78 2.06 8.78 1.22 10.98 1.22
                 10.98 1.86 13.26 1.86 13.26 2.12 13.82 2.12 ;
        RECT  10.90 4.00 13.46 4.32 ;
        POLYGON  12.62 2.92 12.14 2.92 12.14 3.68 9.74 3.68 9.74 3.06 7.64 3.06
                 7.64 2.74 9.74 2.74 9.74 1.86 10.10 1.86 10.10 2.18 10.06 2.18
                 10.06 3.36 11.82 3.36 11.82 2.58 12.62 2.58 ;
        RECT  7.70 3.58 8.90 3.90 ;
        RECT  7.00 1.22 8.46 1.54 ;
        POLYGON  8.46 4.54 6.52 4.54 6.52 4.30 4.14 4.30 4.14 3.70 1.68 3.70
                 1.68 2.42 1.58 2.42 1.58 1.22 1.90 1.22 1.90 2.10 2.00 2.10
                 2.00 3.38 4.46 3.38 4.46 3.98 6.84 3.98 6.84 4.22 8.46 4.22 ;
        POLYGON  7.32 3.70 7.00 3.70 7.00 3.02 5.96 3.02 5.96 2.18 2.96 2.18
                 2.96 2.98 2.64 2.98 2.64 1.86 5.96 1.86 5.96 1.22 6.30 1.22
                 6.30 1.54 6.28 1.54 6.28 2.70 7.32 2.70 ;
        RECT  4.82 3.34 6.62 3.66 ;
        RECT  4.60 1.22 5.60 1.54 ;
        RECT  1.82 4.02 3.63 4.34 ;
        RECT  2.28 1.22 3.28 1.54 ;
        POLYGON  1.36 2.98 1.16 2.98 1.16 3.72 0.50 3.72 0.50 4.54 0.18 4.54
                 0.18 3.40 0.84 3.40 0.84 1.54 0.18 1.54 0.18 1.22 1.16 1.22
                 1.16 2.66 1.36 2.66 ;
    END
END dffprsqb_4

MACRO dffprsqb_2
    CLASS CORE ;
    FOREIGN dffprsqb_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.64 2.72 11.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.72 4.64 3.04 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.96 3.04 20.74 3.04 20.74 4.54 20.42 4.54 20.42 1.22
                 20.74 1.22 20.74 2.72 20.96 2.72 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.12 0.52 3.04 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.28 2.50 3.68 3.06 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 0.90 19.86 0.90 19.86 1.54 19.54 1.54 19.54 0.90
                 16.64 0.90 16.64 1.54 16.32 1.54 16.32 0.90 4.20 0.90
                 4.20 1.54 3.88 1.54 3.88 0.90 0.00 0.90 0.00 -0.90 21.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 6.66 0.00 6.66 0.00 4.86 0.99 4.86 0.99 4.16 1.31 4.16
                 1.31 4.86 5.52 4.86 5.52 4.62 5.84 4.62 5.84 4.86 9.40 4.86
                 9.40 4.16 9.72 4.16 9.72 4.86 11.68 4.86 11.68 4.64 12.00 4.64
                 12.00 4.86 15.32 4.86 15.32 3.94 15.64 3.94 15.64 4.86
                 19.60 4.86 19.60 4.26 19.92 4.26 19.92 4.86 21.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.10 3.06 18.42 3.06 18.42 3.90 18.10 3.90 18.10 3.06
                 17.02 3.06 17.02 4.54 16.70 4.54 16.70 2.86 15.92 2.86
                 15.92 2.54 17.02 2.54 17.02 2.74 18.78 2.74 18.78 1.22
                 19.10 1.22 19.10 2.74 19.78 2.74 19.78 2.62 20.10 2.62 ;
        POLYGON  19.10 4.54 17.40 4.54 17.40 3.58 17.72 3.58 17.72 4.22
                 19.10 4.22 ;
        POLYGON  18.12 2.42 17.79 2.42 17.79 2.18 14.56 2.18 14.56 2.70
                 14.16 3.10 14.16 4.12 13.84 4.12 13.84 2.96 14.24 2.56
                 14.24 1.22 14.56 1.22 14.56 1.86 18.12 1.86 ;
        RECT  17.02 1.22 18.02 1.54 ;
        POLYGON  16.34 3.62 14.86 3.62 14.86 3.80 14.54 3.80 14.54 3.30
                 16.34 3.30 ;
        RECT  14.94 1.22 15.94 1.54 ;
        RECT  11.30 1.22 13.86 1.54 ;
        POLYGON  13.82 2.44 13.26 2.44 13.26 3.68 12.46 3.68 12.46 3.36
                 12.94 3.36 12.94 2.18 10.66 2.18 10.66 1.54 9.10 1.54
                 9.10 2.38 7.04 2.38 7.04 2.06 8.78 2.06 8.78 1.22 10.98 1.22
                 10.98 1.86 13.26 1.86 13.26 2.12 13.82 2.12 ;
        RECT  10.90 4.00 13.46 4.32 ;
        POLYGON  12.62 2.92 12.14 2.92 12.14 3.68 9.74 3.68 9.74 3.06 7.64 3.06
                 7.64 2.74 9.74 2.74 9.74 1.86 10.10 1.86 10.10 2.18 10.06 2.18
                 10.06 3.36 11.82 3.36 11.82 2.58 12.62 2.58 ;
        RECT  7.70 3.58 8.90 3.90 ;
        RECT  7.00 1.22 8.46 1.54 ;
        POLYGON  8.46 4.54 6.52 4.54 6.52 4.30 4.14 4.30 4.14 3.70 1.68 3.70
                 1.68 2.42 1.58 2.42 1.58 1.22 1.90 1.22 1.90 2.10 2.00 2.10
                 2.00 3.38 4.46 3.38 4.46 3.98 6.84 3.98 6.84 4.22 8.46 4.22 ;
        POLYGON  7.32 3.70 7.00 3.70 7.00 3.02 5.96 3.02 5.96 2.18 2.96 2.18
                 2.96 2.98 2.64 2.98 2.64 1.86 5.96 1.86 5.96 1.22 6.30 1.22
                 6.30 1.54 6.28 1.54 6.28 2.70 7.32 2.70 ;
        RECT  4.82 3.34 6.62 3.66 ;
        RECT  4.60 1.22 5.60 1.54 ;
        RECT  1.82 4.02 3.63 4.34 ;
        RECT  2.28 1.22 3.28 1.54 ;
        POLYGON  1.36 2.98 1.16 2.98 1.16 3.72 0.50 3.72 0.50 4.54 0.18 4.54
                 0.18 3.40 0.84 3.40 0.84 1.54 0.18 1.54 0.18 1.22 1.16 1.22
                 1.16 2.66 1.36 2.66 ;
    END
END dffprsqb_2

MACRO dffprsqb_1
    CLASS CORE ;
    FOREIGN dffprsqb_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.64 2.72 11.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.72 4.64 3.04 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.96 3.04 20.74 3.04 20.74 4.54 20.42 4.54 20.42 1.22
                 20.74 1.22 20.74 2.72 20.96 2.72 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.12 0.52 3.04 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.28 2.50 3.68 3.06 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 0.90 19.86 0.90 19.86 1.54 19.54 1.54 19.54 0.90
                 16.64 0.90 16.64 1.54 16.32 1.54 16.32 0.90 4.20 0.90
                 4.20 1.54 3.88 1.54 3.88 0.90 0.00 0.90 0.00 -0.90 21.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 6.66 0.00 6.66 0.00 4.86 0.99 4.86 0.99 4.16 1.31 4.16
                 1.31 4.86 5.52 4.86 5.52 4.62 5.84 4.62 5.84 4.86 9.40 4.86
                 9.40 4.16 9.72 4.16 9.72 4.86 11.68 4.86 11.68 4.64 12.00 4.64
                 12.00 4.86 15.32 4.86 15.32 3.94 15.64 3.94 15.64 4.86
                 19.60 4.86 19.60 4.26 19.92 4.26 19.92 4.86 21.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.10 3.06 18.42 3.06 18.42 3.90 18.10 3.90 18.10 3.06
                 17.02 3.06 17.02 4.54 16.70 4.54 16.70 2.86 15.92 2.86
                 15.92 2.54 17.02 2.54 17.02 2.74 18.78 2.74 18.78 1.22
                 19.10 1.22 19.10 2.74 19.78 2.74 19.78 2.62 20.10 2.62 ;
        POLYGON  19.10 4.54 17.40 4.54 17.40 3.58 17.72 3.58 17.72 4.22
                 19.10 4.22 ;
        POLYGON  18.12 2.42 17.79 2.42 17.79 2.18 14.56 2.18 14.56 2.70
                 14.16 3.10 14.16 4.12 13.84 4.12 13.84 2.96 14.24 2.56
                 14.24 1.22 14.56 1.22 14.56 1.86 18.12 1.86 ;
        RECT  17.02 1.22 18.02 1.54 ;
        POLYGON  16.34 3.62 14.86 3.62 14.86 3.80 14.54 3.80 14.54 3.30
                 16.34 3.30 ;
        RECT  14.94 1.22 15.94 1.54 ;
        RECT  11.30 1.22 13.86 1.54 ;
        POLYGON  13.82 2.44 13.26 2.44 13.26 3.68 12.46 3.68 12.46 3.36
                 12.94 3.36 12.94 2.18 10.66 2.18 10.66 1.54 9.10 1.54
                 9.10 2.38 7.04 2.38 7.04 2.06 8.78 2.06 8.78 1.22 10.98 1.22
                 10.98 1.86 13.26 1.86 13.26 2.12 13.82 2.12 ;
        RECT  10.90 4.00 13.46 4.32 ;
        POLYGON  12.62 2.92 12.14 2.92 12.14 3.68 9.74 3.68 9.74 3.06 7.64 3.06
                 7.64 2.74 9.74 2.74 9.74 1.86 10.10 1.86 10.10 2.18 10.06 2.18
                 10.06 3.36 11.82 3.36 11.82 2.58 12.62 2.58 ;
        RECT  7.70 3.58 8.90 3.90 ;
        RECT  7.00 1.22 8.46 1.54 ;
        POLYGON  8.46 4.54 6.52 4.54 6.52 4.30 4.14 4.30 4.14 3.70 1.68 3.70
                 1.68 2.42 1.58 2.42 1.58 1.22 1.90 1.22 1.90 2.10 2.00 2.10
                 2.00 3.38 4.46 3.38 4.46 3.98 6.84 3.98 6.84 4.22 8.46 4.22 ;
        POLYGON  7.32 3.70 7.00 3.70 7.00 3.02 5.96 3.02 5.96 2.18 2.96 2.18
                 2.96 2.98 2.64 2.98 2.64 1.86 5.96 1.86 5.96 1.22 6.30 1.22
                 6.30 1.54 6.28 1.54 6.28 2.70 7.32 2.70 ;
        RECT  4.82 3.34 6.62 3.66 ;
        RECT  4.60 1.22 5.60 1.54 ;
        RECT  1.82 4.02 3.63 4.34 ;
        RECT  2.28 1.22 3.28 1.54 ;
        POLYGON  1.36 2.98 1.16 2.98 1.16 3.72 0.50 3.72 0.50 4.54 0.18 4.54
                 0.18 3.40 0.84 3.40 0.84 1.54 0.18 1.54 0.18 1.22 1.16 1.22
                 1.16 2.66 1.36 2.66 ;
    END
END dffprsqb_1

MACRO dffprsq_4
    CLASS CORE ;
    FOREIGN dffprsq_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.04 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.64 2.72 11.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.72 4.64 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  22.88 3.04 22.85 3.04 22.85 4.54 22.53 4.54 22.53 3.04
                 21.45 3.04 21.45 4.54 21.13 4.54 21.13 2.75 21.22 2.75
                 21.22 1.55 21.13 1.55 21.13 1.22 21.54 1.22 21.54 2.72
                 22.53 2.72 22.53 1.22 22.85 1.22 22.85 2.72 22.88 2.72 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.12 0.52 3.04 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.28 2.50 3.68 3.06 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  23.04 0.90 19.86 0.90 19.86 1.54 19.54 1.54 19.54 0.90
                 16.64 0.90 16.64 1.54 16.32 1.54 16.32 0.90 4.20 0.90
                 4.20 1.54 3.88 1.54 3.88 0.90 0.00 0.90 0.00 -0.90 23.04 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  23.04 6.66 0.00 6.66 0.00 4.86 0.99 4.86 0.99 4.16 1.31 4.16
                 1.31 4.86 5.52 4.86 5.52 4.62 5.84 4.62 5.84 4.86 9.40 4.86
                 9.40 4.16 9.72 4.16 9.72 4.86 11.68 4.86 11.68 4.64 12.00 4.64
                 12.00 4.86 15.32 4.86 15.32 3.94 15.64 3.94 15.64 4.86
                 19.60 4.86 19.60 4.22 19.92 4.22 19.92 4.86 21.83 4.86
                 21.83 3.58 22.15 3.58 22.15 4.86 23.04 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.90 2.52 20.74 2.52 20.74 4.54 20.42 4.54 20.42 1.22
                 20.74 1.22 20.74 2.20 20.90 2.20 ;
        POLYGON  20.10 3.06 18.42 3.06 18.42 3.90 18.10 3.90 18.10 3.06
                 17.02 3.06 17.02 4.54 16.70 4.54 16.70 2.86 15.92 2.86
                 15.92 2.54 17.02 2.54 17.02 2.74 18.78 2.74 18.78 1.22
                 19.10 1.22 19.10 2.74 19.78 2.74 19.78 2.62 20.10 2.62 ;
        POLYGON  19.10 4.54 17.40 4.54 17.40 3.58 17.72 3.58 17.72 4.22
                 19.10 4.22 ;
        POLYGON  18.12 2.42 17.79 2.42 17.79 2.18 14.56 2.18 14.56 2.70
                 14.16 3.10 14.16 4.12 13.84 4.12 13.84 2.96 14.24 2.56
                 14.24 1.22 14.56 1.22 14.56 1.86 18.12 1.86 ;
        RECT  17.02 1.22 18.02 1.54 ;
        POLYGON  16.34 3.62 14.86 3.62 14.86 3.80 14.54 3.80 14.54 3.30
                 16.34 3.30 ;
        RECT  14.94 1.22 15.94 1.54 ;
        RECT  11.30 1.22 13.86 1.54 ;
        POLYGON  13.82 2.44 13.26 2.44 13.26 3.68 12.46 3.68 12.46 3.36
                 12.94 3.36 12.94 2.18 10.66 2.18 10.66 1.54 9.10 1.54
                 9.10 2.38 7.04 2.38 7.04 2.06 8.78 2.06 8.78 1.22 10.98 1.22
                 10.98 1.86 13.26 1.86 13.26 2.12 13.82 2.12 ;
        RECT  10.90 4.00 13.46 4.32 ;
        POLYGON  12.62 2.92 12.14 2.92 12.14 3.68 9.74 3.68 9.74 3.06 7.64 3.06
                 7.64 2.74 9.74 2.74 9.74 1.86 10.10 1.86 10.10 2.18 10.06 2.18
                 10.06 3.36 11.82 3.36 11.82 2.58 12.62 2.58 ;
        RECT  7.70 3.58 8.90 3.90 ;
        RECT  7.00 1.22 8.46 1.54 ;
        POLYGON  8.46 4.54 6.52 4.54 6.52 4.30 4.14 4.30 4.14 3.70 1.68 3.70
                 1.68 2.42 1.58 2.42 1.58 1.22 1.90 1.22 1.90 2.10 2.00 2.10
                 2.00 3.38 4.46 3.38 4.46 3.98 6.84 3.98 6.84 4.22 8.46 4.22 ;
        POLYGON  7.32 3.70 7.00 3.70 7.00 3.02 5.96 3.02 5.96 2.18 2.96 2.18
                 2.96 2.98 2.64 2.98 2.64 1.86 5.96 1.86 5.96 1.22 6.30 1.22
                 6.30 1.54 6.28 1.54 6.28 2.70 7.32 2.70 ;
        RECT  4.82 3.34 6.62 3.66 ;
        RECT  4.60 1.22 5.60 1.54 ;
        RECT  1.82 4.02 3.63 4.34 ;
        RECT  2.28 1.22 3.28 1.54 ;
        POLYGON  1.36 2.98 1.16 2.98 1.16 3.72 0.50 3.72 0.50 4.54 0.18 4.54
                 0.18 3.40 0.84 3.40 0.84 1.54 0.18 1.54 0.18 1.22 1.16 1.22
                 1.16 2.66 1.36 2.66 ;
    END
END dffprsq_4

MACRO dffprsq_2
    CLASS CORE ;
    FOREIGN dffprsq_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.64 2.72 11.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.72 4.64 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  22.24 3.04 22.12 3.04 22.12 4.54 21.80 4.54 21.80 1.64
                 22.12 1.64 22.12 2.72 22.24 2.72 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.12 0.52 3.04 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.28 2.50 3.68 3.06 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  22.40 0.90 21.42 0.90 21.42 1.48 21.10 1.48 21.10 0.90
                 19.86 0.90 19.86 1.54 19.54 1.54 19.54 0.90 16.64 0.90
                 16.64 1.54 16.32 1.54 16.32 0.90 4.20 0.90 4.20 1.54 3.88 1.54
                 3.88 0.90 0.00 0.90 0.00 -0.90 22.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  22.40 6.66 0.00 6.66 0.00 4.86 0.99 4.86 0.99 4.16 1.31 4.16
                 1.31 4.86 5.52 4.86 5.52 4.62 5.84 4.62 5.84 4.86 9.40 4.86
                 9.40 4.16 9.72 4.16 9.72 4.86 11.68 4.86 11.68 4.64 12.00 4.64
                 12.00 4.86 15.32 4.86 15.32 3.94 15.64 3.94 15.64 4.86
                 19.60 4.86 19.60 4.26 19.92 4.26 19.92 4.86 21.10 4.86
                 21.10 4.22 21.42 4.22 21.42 4.86 22.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.92 2.86 20.74 2.86 20.74 4.54 20.42 4.54 20.42 1.22
                 20.74 1.22 20.74 2.54 20.92 2.54 ;
        POLYGON  20.10 3.06 18.42 3.06 18.42 3.90 18.10 3.90 18.10 3.06
                 17.02 3.06 17.02 4.54 16.70 4.54 16.70 2.86 15.92 2.86
                 15.92 2.54 17.02 2.54 17.02 2.74 18.78 2.74 18.78 1.22
                 19.10 1.22 19.10 2.74 19.78 2.74 19.78 2.62 20.10 2.62 ;
        POLYGON  19.10 4.54 17.40 4.54 17.40 3.58 17.72 3.58 17.72 4.22
                 19.10 4.22 ;
        POLYGON  18.12 2.42 17.79 2.42 17.79 2.18 14.56 2.18 14.56 2.70
                 14.16 3.10 14.16 4.12 13.84 4.12 13.84 2.96 14.24 2.56
                 14.24 1.22 14.56 1.22 14.56 1.86 18.12 1.86 ;
        RECT  17.02 1.22 18.02 1.54 ;
        POLYGON  16.34 3.62 14.86 3.62 14.86 3.80 14.54 3.80 14.54 3.30
                 16.34 3.30 ;
        RECT  14.94 1.22 15.94 1.54 ;
        RECT  11.30 1.22 13.86 1.54 ;
        POLYGON  13.82 2.44 13.26 2.44 13.26 3.68 12.46 3.68 12.46 3.36
                 12.94 3.36 12.94 2.18 10.66 2.18 10.66 1.54 9.10 1.54
                 9.10 2.38 7.04 2.38 7.04 2.06 8.78 2.06 8.78 1.22 10.98 1.22
                 10.98 1.86 13.26 1.86 13.26 2.12 13.82 2.12 ;
        RECT  10.90 4.00 13.46 4.32 ;
        POLYGON  12.62 2.92 12.14 2.92 12.14 3.68 9.74 3.68 9.74 3.06 7.64 3.06
                 7.64 2.74 9.74 2.74 9.74 1.86 10.10 1.86 10.10 2.18 10.06 2.18
                 10.06 3.36 11.82 3.36 11.82 2.58 12.62 2.58 ;
        RECT  7.70 3.58 8.90 3.90 ;
        RECT  7.00 1.22 8.46 1.54 ;
        POLYGON  8.46 4.54 6.52 4.54 6.52 4.30 4.14 4.30 4.14 3.70 1.68 3.70
                 1.68 2.42 1.58 2.42 1.58 1.22 1.90 1.22 1.90 2.10 2.00 2.10
                 2.00 3.38 4.46 3.38 4.46 3.98 6.84 3.98 6.84 4.22 8.46 4.22 ;
        POLYGON  7.32 3.70 7.00 3.70 7.00 3.02 5.96 3.02 5.96 2.18 2.96 2.18
                 2.96 2.98 2.64 2.98 2.64 1.86 5.96 1.86 5.96 1.22 6.30 1.22
                 6.30 1.54 6.28 1.54 6.28 2.70 7.32 2.70 ;
        RECT  4.82 3.34 6.62 3.66 ;
        RECT  4.60 1.22 5.60 1.54 ;
        RECT  1.82 4.02 3.63 4.34 ;
        RECT  2.28 1.22 3.28 1.54 ;
        POLYGON  1.36 2.98 1.16 2.98 1.16 3.72 0.50 3.72 0.50 4.54 0.18 4.54
                 0.18 3.40 0.84 3.40 0.84 1.54 0.18 1.54 0.18 1.22 1.16 1.22
                 1.16 2.66 1.36 2.66 ;
    END
END dffprsq_2

MACRO dffprsq_1
    CLASS CORE ;
    FOREIGN dffprsq_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.64 2.72 11.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.72 4.64 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  22.24 3.04 22.12 3.04 22.12 4.54 21.80 4.54 21.80 1.22
                 22.12 1.22 22.12 2.72 22.24 2.72 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.12 0.52 3.04 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.28 2.50 3.68 3.06 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  22.40 0.90 21.42 0.90 21.42 1.54 21.10 1.54 21.10 0.90
                 19.86 0.90 19.86 1.54 19.54 1.54 19.54 0.90 16.64 0.90
                 16.64 1.54 16.32 1.54 16.32 0.90 4.20 0.90 4.20 1.54 3.88 1.54
                 3.88 0.90 0.00 0.90 0.00 -0.90 22.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  22.40 6.66 0.00 6.66 0.00 4.86 0.99 4.86 0.99 4.16 1.31 4.16
                 1.31 4.86 5.52 4.86 5.52 4.62 5.84 4.62 5.84 4.86 9.40 4.86
                 9.40 4.16 9.72 4.16 9.72 4.86 11.68 4.86 11.68 4.64 12.00 4.64
                 12.00 4.86 15.32 4.86 15.32 3.94 15.64 3.94 15.64 4.86
                 19.60 4.86 19.60 4.28 19.92 4.28 19.92 4.86 21.10 4.86
                 21.10 4.28 21.42 4.28 21.42 4.86 22.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.92 2.86 20.74 2.86 20.74 4.54 20.42 4.54 20.42 1.22
                 20.74 1.22 20.74 2.54 20.92 2.54 ;
        POLYGON  20.10 3.06 18.42 3.06 18.42 3.90 18.10 3.90 18.10 3.06
                 17.02 3.06 17.02 4.54 16.70 4.54 16.70 2.86 15.92 2.86
                 15.92 2.54 17.02 2.54 17.02 2.74 18.78 2.74 18.78 1.22
                 19.10 1.22 19.10 2.74 19.78 2.74 19.78 2.62 20.10 2.62 ;
        POLYGON  19.10 4.54 17.40 4.54 17.40 3.58 17.72 3.58 17.72 4.22
                 19.10 4.22 ;
        POLYGON  18.12 2.42 17.79 2.42 17.79 2.18 14.56 2.18 14.56 2.70
                 14.16 3.10 14.16 4.12 13.84 4.12 13.84 2.96 14.24 2.56
                 14.24 1.22 14.56 1.22 14.56 1.86 18.12 1.86 ;
        RECT  17.02 1.22 18.02 1.54 ;
        POLYGON  16.34 3.62 14.86 3.62 14.86 3.80 14.54 3.80 14.54 3.30
                 16.34 3.30 ;
        RECT  14.94 1.22 15.94 1.54 ;
        RECT  11.30 1.22 13.86 1.54 ;
        POLYGON  13.82 2.44 13.26 2.44 13.26 3.68 12.46 3.68 12.46 3.36
                 12.94 3.36 12.94 2.18 10.66 2.18 10.66 1.54 9.10 1.54
                 9.10 2.38 7.04 2.38 7.04 2.06 8.78 2.06 8.78 1.22 10.98 1.22
                 10.98 1.86 13.26 1.86 13.26 2.12 13.82 2.12 ;
        RECT  10.90 4.00 13.46 4.32 ;
        POLYGON  12.62 2.92 12.14 2.92 12.14 3.68 9.74 3.68 9.74 3.06 7.64 3.06
                 7.64 2.74 9.74 2.74 9.74 1.86 10.10 1.86 10.10 2.18 10.06 2.18
                 10.06 3.36 11.82 3.36 11.82 2.58 12.62 2.58 ;
        RECT  7.70 3.58 8.90 3.90 ;
        RECT  7.00 1.22 8.46 1.54 ;
        POLYGON  8.46 4.54 6.52 4.54 6.52 4.30 4.14 4.30 4.14 3.70 1.68 3.70
                 1.68 2.42 1.58 2.42 1.58 1.22 1.90 1.22 1.90 2.10 2.00 2.10
                 2.00 3.38 4.46 3.38 4.46 3.98 6.84 3.98 6.84 4.22 8.46 4.22 ;
        POLYGON  7.32 3.70 7.00 3.70 7.00 3.02 5.96 3.02 5.96 2.18 2.96 2.18
                 2.96 2.98 2.64 2.98 2.64 1.86 5.96 1.86 5.96 1.22 6.30 1.22
                 6.30 1.54 6.28 1.54 6.28 2.70 7.32 2.70 ;
        RECT  4.82 3.34 6.62 3.66 ;
        RECT  4.60 1.22 5.60 1.54 ;
        RECT  1.82 4.02 3.63 4.34 ;
        RECT  2.28 1.22 3.28 1.54 ;
        POLYGON  1.36 2.98 1.16 2.98 1.16 3.72 0.50 3.72 0.50 4.54 0.18 4.54
                 0.18 3.40 0.84 3.40 0.84 1.54 0.18 1.54 0.18 1.22 1.16 1.22
                 1.16 2.66 1.36 2.66 ;
    END
END dffprsq_1

MACRO dffprs_4
    CLASS CORE ;
    FOREIGN dffprs_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 25.60 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.64 2.72 11.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.72 4.64 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  23.52 3.25 21.58 3.25 21.58 2.93 23.20 2.93 23.20 2.52
                 22.97 2.52 22.97 1.54 21.10 1.54 21.10 1.22 23.29 1.22
                 23.29 2.20 23.52 2.20 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  25.44 4.53 23.67 4.53 23.67 4.21 25.12 4.21 25.12 1.90
                 23.67 1.90 23.67 1.58 25.44 1.58 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.12 0.52 3.04 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.28 2.50 3.68 3.06 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  25.60 0.90 19.86 0.90 19.86 1.54 19.54 1.54 19.54 0.90
                 16.64 0.90 16.64 1.54 16.32 1.54 16.32 0.90 4.20 0.90
                 4.20 1.54 3.88 1.54 3.88 0.90 0.00 0.90 0.00 -0.90 25.60 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  25.60 6.66 0.00 6.66 0.00 4.86 0.99 4.86 0.99 4.16 1.31 4.16
                 1.31 4.86 5.52 4.86 5.52 4.62 5.84 4.62 5.84 4.86 9.40 4.86
                 9.40 4.16 9.72 4.16 9.72 4.86 11.68 4.86 11.68 4.64 12.00 4.64
                 12.00 4.86 15.32 4.86 15.32 3.94 15.64 3.94 15.64 4.86
                 19.60 4.86 19.60 4.64 19.92 4.64 19.92 4.86 22.24 4.86
                 22.24 4.81 22.64 4.81 22.64 4.86 25.60 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  24.69 3.89 22.03 3.89 22.03 4.18 19.78 4.18 19.78 3.06
                 18.42 3.06 18.42 3.90 18.10 3.90 18.10 3.06 17.02 3.06
                 17.02 4.54 16.70 4.54 16.70 2.86 15.92 2.86 15.92 2.54
                 17.02 2.54 17.02 2.74 18.78 2.74 18.78 1.22 19.10 1.22
                 19.10 2.74 19.78 2.74 19.78 2.62 20.10 2.62 20.10 3.86
                 21.71 3.86 21.71 3.57 24.37 3.57 24.37 2.34 24.69 2.34 ;
        POLYGON  20.92 2.55 20.74 2.55 20.74 3.42 20.42 3.42 20.42 1.22
                 20.74 1.22 20.74 2.23 20.92 2.23 ;
        POLYGON  19.10 4.54 17.40 4.54 17.40 3.58 17.72 3.58 17.72 4.22
                 19.10 4.22 ;
        POLYGON  18.12 2.42 17.79 2.42 17.79 2.18 14.56 2.18 14.56 2.70
                 14.16 3.10 14.16 4.12 13.84 4.12 13.84 2.96 14.24 2.56
                 14.24 1.22 14.56 1.22 14.56 1.86 18.12 1.86 ;
        RECT  17.02 1.22 18.02 1.54 ;
        POLYGON  16.34 3.62 14.86 3.62 14.86 3.80 14.54 3.80 14.54 3.30
                 16.34 3.30 ;
        RECT  14.94 1.22 15.94 1.54 ;
        RECT  11.30 1.22 13.86 1.54 ;
        POLYGON  13.82 2.44 13.26 2.44 13.26 3.68 12.46 3.68 12.46 3.36
                 12.94 3.36 12.94 2.18 10.66 2.18 10.66 1.54 9.10 1.54
                 9.10 2.38 7.04 2.38 7.04 2.06 8.78 2.06 8.78 1.22 10.98 1.22
                 10.98 1.86 13.26 1.86 13.26 2.12 13.82 2.12 ;
        RECT  10.90 4.00 13.46 4.32 ;
        POLYGON  12.62 2.92 12.14 2.92 12.14 3.68 9.74 3.68 9.74 3.06 7.64 3.06
                 7.64 2.74 9.74 2.74 9.74 1.86 10.10 1.86 10.10 2.18 10.06 2.18
                 10.06 3.36 11.82 3.36 11.82 2.58 12.62 2.58 ;
        RECT  7.70 3.58 8.90 3.90 ;
        RECT  7.00 1.22 8.46 1.54 ;
        POLYGON  8.46 4.54 6.52 4.54 6.52 4.30 4.14 4.30 4.14 3.70 1.68 3.70
                 1.68 2.42 1.58 2.42 1.58 1.22 1.90 1.22 1.90 2.10 2.00 2.10
                 2.00 3.38 4.46 3.38 4.46 3.98 6.84 3.98 6.84 4.22 8.46 4.22 ;
        POLYGON  7.32 3.70 7.00 3.70 7.00 3.02 5.96 3.02 5.96 2.18 2.96 2.18
                 2.96 2.98 2.64 2.98 2.64 1.86 5.96 1.86 5.96 1.22 6.30 1.22
                 6.30 1.54 6.28 1.54 6.28 2.70 7.32 2.70 ;
        RECT  4.82 3.34 6.62 3.66 ;
        RECT  4.60 1.22 5.60 1.54 ;
        RECT  1.82 4.02 3.63 4.34 ;
        RECT  2.28 1.22 3.28 1.54 ;
        POLYGON  1.36 2.98 1.16 2.98 1.16 3.72 0.50 3.72 0.50 4.54 0.18 4.54
                 0.18 3.40 0.84 3.40 0.84 1.54 0.18 1.54 0.18 1.22 1.16 1.22
                 1.16 2.66 1.36 2.66 ;
    END
END dffprs_4

MACRO dffprs_2
    CLASS CORE ;
    FOREIGN dffprs_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.04 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.64 2.72 11.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.72 4.64 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  21.60 3.45 21.10 3.45 21.10 3.13 21.28 3.13 21.28 2.27
                 21.10 2.27 21.10 1.22 21.42 1.22 21.42 1.95 21.60 1.95 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  22.88 4.54 22.54 4.54 22.54 4.22 22.56 4.22 22.56 1.54
                 22.54 1.54 22.54 1.22 22.88 1.22 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.12 0.52 3.04 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.28 2.50 3.68 3.06 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  23.04 0.90 22.12 0.90 22.12 1.54 21.80 1.54 21.80 0.90
                 19.86 0.90 19.86 1.54 19.54 1.54 19.54 0.90 16.64 0.90
                 16.64 1.54 16.32 1.54 16.32 0.90 4.20 0.90 4.20 1.54 3.88 1.54
                 3.88 0.90 0.00 0.90 0.00 -0.90 23.04 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  23.04 6.66 0.00 6.66 0.00 4.86 0.99 4.86 0.99 4.16 1.31 4.16
                 1.31 4.86 5.52 4.86 5.52 4.62 5.84 4.62 5.84 4.86 9.40 4.86
                 9.40 4.16 9.72 4.16 9.72 4.86 11.68 4.86 11.68 4.64 12.00 4.64
                 12.00 4.86 15.32 4.86 15.32 3.94 15.64 3.94 15.64 4.86
                 19.60 4.86 19.60 4.41 19.92 4.41 19.92 4.86 23.04 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  22.24 4.09 19.78 4.09 19.78 3.06 18.42 3.06 18.42 3.90
                 18.10 3.90 18.10 3.06 17.02 3.06 17.02 4.54 16.70 4.54
                 16.70 2.86 15.92 2.86 15.92 2.54 17.02 2.54 17.02 2.74
                 18.78 2.74 18.78 1.22 19.10 1.22 19.10 2.74 19.78 2.74
                 19.78 2.62 20.10 2.62 20.10 3.77 21.92 3.77 21.92 2.38
                 22.24 2.38 ;
        POLYGON  20.92 2.86 20.74 2.86 20.74 3.42 20.42 3.42 20.42 1.22
                 20.74 1.22 20.74 2.54 20.92 2.54 ;
        POLYGON  19.10 4.54 17.40 4.54 17.40 3.58 17.72 3.58 17.72 4.22
                 18.78 4.22 18.78 3.58 19.10 3.58 ;
        POLYGON  18.12 2.42 17.79 2.42 17.79 2.18 14.56 2.18 14.56 2.70
                 14.16 3.10 14.16 4.12 13.84 4.12 13.84 2.96 14.24 2.56
                 14.24 1.22 14.56 1.22 14.56 1.86 18.12 1.86 ;
        RECT  17.02 1.22 18.02 1.54 ;
        POLYGON  16.34 3.62 14.86 3.62 14.86 3.80 14.54 3.80 14.54 3.30
                 16.34 3.30 ;
        RECT  14.94 1.22 15.94 1.54 ;
        RECT  11.30 1.22 13.86 1.54 ;
        POLYGON  13.82 2.44 13.26 2.44 13.26 3.68 12.46 3.68 12.46 3.36
                 12.94 3.36 12.94 2.18 10.66 2.18 10.66 1.54 9.10 1.54
                 9.10 2.38 7.04 2.38 7.04 2.06 8.78 2.06 8.78 1.22 10.98 1.22
                 10.98 1.86 13.26 1.86 13.26 2.12 13.82 2.12 ;
        RECT  10.90 4.00 13.46 4.32 ;
        POLYGON  12.62 2.92 12.14 2.92 12.14 3.68 9.74 3.68 9.74 3.06 7.64 3.06
                 7.64 2.74 9.74 2.74 9.74 1.86 10.10 1.86 10.10 2.18 10.06 2.18
                 10.06 3.36 11.82 3.36 11.82 2.58 12.62 2.58 ;
        RECT  7.70 3.58 8.90 3.90 ;
        RECT  7.00 1.22 8.46 1.54 ;
        POLYGON  8.46 4.54 6.52 4.54 6.52 4.30 4.14 4.30 4.14 3.70 1.68 3.70
                 1.68 2.42 1.58 2.42 1.58 1.22 1.90 1.22 1.90 2.10 2.00 2.10
                 2.00 3.38 4.46 3.38 4.46 3.98 6.84 3.98 6.84 4.22 8.46 4.22 ;
        POLYGON  7.32 3.70 7.00 3.70 7.00 3.02 5.96 3.02 5.96 2.18 2.96 2.18
                 2.96 2.98 2.64 2.98 2.64 1.86 5.96 1.86 5.96 1.22 6.30 1.22
                 6.30 1.54 6.28 1.54 6.28 2.70 7.32 2.70 ;
        RECT  4.82 3.34 6.62 3.66 ;
        RECT  4.60 1.22 5.60 1.54 ;
        RECT  1.82 4.02 3.63 4.34 ;
        RECT  2.28 1.22 3.28 1.54 ;
        POLYGON  1.36 2.98 1.16 2.98 1.16 3.72 0.50 3.72 0.50 4.54 0.18 4.54
                 0.18 3.40 0.84 3.40 0.84 1.54 0.18 1.54 0.18 1.22 1.16 1.22
                 1.16 2.66 1.36 2.66 ;
    END
END dffprs_2

MACRO dffprs_1
    CLASS CORE ;
    FOREIGN dffprs_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.04 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.64 2.72 11.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.72 4.64 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.21  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  21.60 3.45 21.10 3.45 21.10 3.13 21.28 3.13 21.28 2.27
                 21.10 2.27 21.10 1.22 21.42 1.22 21.42 1.95 21.60 1.95 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.21  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  22.88 4.54 22.54 4.54 22.54 4.22 22.56 4.22 22.56 1.54
                 22.54 1.54 22.54 1.22 22.88 1.22 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.12 0.52 3.04 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.28 2.50 3.68 3.06 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  23.04 0.90 22.12 0.90 22.12 1.54 21.80 1.54 21.80 0.90
                 19.86 0.90 19.86 1.54 19.54 1.54 19.54 0.90 16.64 0.90
                 16.64 1.54 16.32 1.54 16.32 0.90 4.20 0.90 4.20 1.54 3.88 1.54
                 3.88 0.90 0.00 0.90 0.00 -0.90 23.04 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  23.04 6.66 0.00 6.66 0.00 4.86 0.99 4.86 0.99 4.16 1.31 4.16
                 1.31 4.86 5.52 4.86 5.52 4.62 5.84 4.62 5.84 4.86 9.40 4.86
                 9.40 4.16 9.72 4.16 9.72 4.86 11.68 4.86 11.68 4.64 12.00 4.64
                 12.00 4.86 15.32 4.86 15.32 3.94 15.64 3.94 15.64 4.86
                 19.66 4.86 19.66 4.41 19.98 4.41 19.98 4.86 21.80 4.86
                 21.80 4.41 22.12 4.41 22.12 4.86 23.04 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  22.24 4.09 19.78 4.09 19.78 3.06 18.42 3.06 18.42 3.90
                 18.10 3.90 18.10 3.06 17.02 3.06 17.02 4.54 16.70 4.54
                 16.70 2.86 15.92 2.86 15.92 2.54 17.02 2.54 17.02 2.74
                 18.78 2.74 18.78 1.22 19.10 1.22 19.10 2.74 19.78 2.74
                 19.78 2.62 20.10 2.62 20.10 3.77 21.92 3.77 21.92 2.38
                 22.24 2.38 ;
        POLYGON  20.92 2.86 20.74 2.86 20.74 3.42 20.42 3.42 20.42 1.22
                 20.74 1.22 20.74 2.54 20.92 2.54 ;
        POLYGON  19.10 4.54 17.40 4.54 17.40 3.58 17.72 3.58 17.72 4.22
                 18.78 4.22 18.78 3.58 19.10 3.58 ;
        POLYGON  18.12 2.42 17.79 2.42 17.79 2.18 14.56 2.18 14.56 2.70
                 14.16 3.10 14.16 4.12 13.84 4.12 13.84 2.96 14.24 2.56
                 14.24 1.22 14.56 1.22 14.56 1.86 18.12 1.86 ;
        RECT  17.02 1.22 18.02 1.54 ;
        POLYGON  16.34 3.62 14.86 3.62 14.86 3.80 14.54 3.80 14.54 3.30
                 16.34 3.30 ;
        RECT  14.94 1.22 15.94 1.54 ;
        RECT  11.30 1.22 13.86 1.54 ;
        POLYGON  13.82 2.44 13.26 2.44 13.26 3.68 12.46 3.68 12.46 3.36
                 12.94 3.36 12.94 2.18 10.66 2.18 10.66 1.54 9.10 1.54
                 9.10 2.38 7.04 2.38 7.04 2.06 8.78 2.06 8.78 1.22 10.98 1.22
                 10.98 1.86 13.26 1.86 13.26 2.12 13.82 2.12 ;
        RECT  10.90 4.00 13.46 4.32 ;
        POLYGON  12.62 2.92 12.14 2.92 12.14 3.68 9.74 3.68 9.74 3.06 7.64 3.06
                 7.64 2.74 9.74 2.74 9.74 1.86 10.10 1.86 10.10 2.18 10.06 2.18
                 10.06 3.36 11.82 3.36 11.82 2.58 12.62 2.58 ;
        RECT  7.70 3.58 8.90 3.90 ;
        RECT  7.00 1.22 8.46 1.54 ;
        POLYGON  8.46 4.54 6.52 4.54 6.52 4.30 4.14 4.30 4.14 3.70 1.68 3.70
                 1.68 2.42 1.58 2.42 1.58 1.22 1.90 1.22 1.90 2.10 2.00 2.10
                 2.00 3.38 4.46 3.38 4.46 3.98 6.84 3.98 6.84 4.22 8.46 4.22 ;
        POLYGON  7.32 3.70 7.00 3.70 7.00 3.02 5.96 3.02 5.96 2.18 2.96 2.18
                 2.96 2.98 2.64 2.98 2.64 1.86 5.96 1.86 5.96 1.22 6.30 1.22
                 6.30 1.54 6.28 1.54 6.28 2.70 7.32 2.70 ;
        RECT  4.82 3.34 6.62 3.66 ;
        RECT  4.60 1.22 5.60 1.54 ;
        RECT  1.82 4.02 3.63 4.34 ;
        RECT  2.28 1.22 3.28 1.54 ;
        POLYGON  1.36 2.98 1.16 2.98 1.16 3.72 0.50 3.72 0.50 4.54 0.18 4.54
                 0.18 3.40 0.84 3.40 0.84 1.54 0.18 1.54 0.18 1.22 1.16 1.22
                 1.16 2.66 1.36 2.66 ;
    END
END dffprs_1

MACRO dffprqb_4
    CLASS CORE ;
    FOREIGN dffprqb_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  7.84 2.72 8.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.08 3.04 2.44 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.96 4.53 19.08 4.53 19.08 4.21 20.64 4.21 20.64 1.90
                 19.08 1.90 19.08 1.58 20.96 1.58 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.22  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 2.08 2.44 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 0.90 20.10 0.90 20.10 1.23 19.78 1.23 19.78 0.90
                 17.78 0.90 17.78 1.54 17.46 1.54 17.46 0.90 8.36 0.90
                 8.36 1.54 8.04 1.54 8.04 0.90 1.20 0.90 1.20 1.54 0.88 1.54
                 0.88 0.90 0.00 0.90 0.00 -0.90 21.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 6.66 0.00 6.66 0.00 4.86 16.08 4.86 16.08 4.20
                 16.40 4.20 16.40 4.86 17.58 4.86 17.58 4.56 17.90 4.56
                 17.90 4.86 21.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.10 3.89 18.72 3.89 18.72 4.54 18.40 4.54 18.40 3.22
                 16.14 3.22 16.14 2.90 18.28 2.90 18.28 2.02 18.16 2.02
                 18.16 1.22 18.48 1.22 18.48 1.76 18.60 1.76 18.60 2.90
                 18.72 2.90 18.72 3.57 19.78 3.57 19.78 2.65 19.74 2.65
                 19.74 2.33 20.10 2.33 ;
        POLYGON  17.94 2.58 15.82 2.58 15.82 3.54 17.08 3.54 17.08 4.54
                 16.76 4.54 16.76 3.86 14.40 3.86 14.22 4.04 14.22 4.54
                 13.90 4.54 13.90 3.90 14.26 3.54 15.50 3.54 15.50 2.58
                 14.82 2.58 14.00 1.76 14.00 1.22 14.32 1.22 14.32 1.62
                 14.96 2.26 17.94 2.26 ;
        RECT  16.08 1.22 17.08 1.54 ;
        RECT  14.70 1.22 15.70 1.54 ;
        RECT  14.60 4.20 15.70 4.52 ;
        POLYGON  14.06 2.60 13.74 2.60 13.74 3.24 13.08 3.90 11.98 3.90
                 11.98 4.54 8.18 4.54 8.18 4.05 8.03 3.90 6.86 3.90 6.86 3.26
                 5.90 3.26 5.90 2.94 7.18 2.94 7.18 3.58 8.17 3.58 8.50 3.91
                 8.50 4.22 11.66 4.22 11.66 3.58 12.94 3.58 13.42 3.10
                 13.42 2.50 13.10 2.18 10.38 2.18 10.38 1.86 13.24 1.86
                 13.66 2.28 14.06 2.28 ;
        RECT  12.62 1.22 13.62 1.54 ;
        RECT  12.52 4.22 13.52 4.54 ;
        POLYGON  13.10 2.96 11.34 2.96 11.34 3.90 8.82 3.90 8.82 2.18 5.58 2.18
                 5.58 3.26 5.26 3.26 5.26 1.86 9.14 1.86 9.14 3.58 11.02 3.58
                 11.02 2.64 13.10 2.64 ;
        POLYGON  12.24 1.54 10.06 1.54 10.06 2.54 10.60 2.54 10.60 2.86
                 9.74 2.86 9.74 1.22 12.24 1.22 ;
        POLYGON  7.86 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 7.86 4.22 ;
        RECT  6.66 1.22 7.66 1.54 ;
        RECT  5.54 3.58 6.54 3.90 ;
        RECT  5.28 1.22 6.28 1.54 ;
        POLYGON  5.08 3.90 4.62 3.90 4.62 2.40 3.68 2.40 3.68 3.08 2.14 3.08
                 2.14 3.90 1.82 3.90 1.82 3.08 0.80 3.08 0.80 2.72 1.12 2.72
                 1.12 2.76 3.36 2.76 3.36 2.08 4.58 2.08 4.58 1.22 4.90 1.22
                 4.90 2.08 4.94 2.08 4.94 3.58 5.08 3.58 ;
        POLYGON  4.30 3.90 2.50 3.90 2.50 3.58 3.98 3.58 3.98 3.36 4.30 3.36 ;
        RECT  3.20 1.22 4.20 1.54 ;
        RECT  1.58 1.22 2.82 1.54 ;
    END
END dffprqb_4

MACRO dffprqb_2
    CLASS CORE ;
    FOREIGN dffprqb_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 20.48 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  7.84 2.72 8.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.08 3.04 2.44 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.19  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.32 4.54 19.92 4.54 19.92 4.22 20.00 4.22 20.00 1.58
                 19.92 1.58 19.92 1.26 20.32 1.26 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.22  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 2.08 2.44 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 0.90 19.40 0.90 19.40 1.58 19.08 1.58 19.08 0.90
                 17.78 0.90 17.78 1.54 17.46 1.54 17.46 0.90 8.36 0.90
                 8.36 1.54 8.04 1.54 8.04 0.90 1.20 0.90 1.20 1.54 0.88 1.54
                 0.88 0.90 0.00 0.90 0.00 -0.90 20.48 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 6.66 0.00 6.66 0.00 4.86 16.08 4.86 16.08 4.12
                 16.40 4.12 16.40 4.86 17.58 4.86 17.58 4.56 17.90 4.56
                 17.90 4.86 20.48 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  19.62 3.91 19.25 4.28 18.28 4.28 18.28 3.16 16.14 3.16
                 16.14 2.84 18.28 2.84 18.28 1.54 18.16 1.54 18.16 1.22
                 18.60 1.22 18.60 3.96 19.09 3.96 19.30 3.75 19.30 2.46
                 19.26 2.46 19.26 2.14 19.62 2.14 ;
        POLYGON  17.96 2.52 15.82 2.52 15.82 3.48 17.08 3.48 17.08 4.54
                 16.76 4.54 16.76 3.80 14.46 3.80 14.22 4.04 14.22 4.54
                 13.90 4.54 13.90 3.90 14.32 3.48 15.50 3.48 15.50 2.52
                 14.76 2.52 14.00 1.76 14.00 1.22 14.32 1.22 14.32 1.62
                 14.90 2.20 17.96 2.20 ;
        RECT  16.08 1.22 17.08 1.54 ;
        RECT  14.70 1.22 15.70 1.54 ;
        RECT  14.60 4.12 15.70 4.44 ;
        POLYGON  14.06 2.60 13.74 2.60 13.74 3.24 13.08 3.90 11.98 3.90
                 11.98 4.54 8.18 4.54 8.18 4.05 8.03 3.90 6.86 3.90 6.86 3.26
                 5.90 3.26 5.90 2.94 7.18 2.94 7.18 3.58 8.17 3.58 8.50 3.91
                 8.50 4.22 11.66 4.22 11.66 3.58 12.94 3.58 13.42 3.10
                 13.42 2.50 13.10 2.18 10.38 2.18 10.38 1.86 13.24 1.86
                 13.66 2.28 14.06 2.28 ;
        RECT  12.62 1.22 13.62 1.54 ;
        RECT  12.52 4.22 13.52 4.54 ;
        POLYGON  13.10 2.96 11.34 2.96 11.34 3.90 8.82 3.90 8.82 2.18 5.58 2.18
                 5.58 3.26 5.26 3.26 5.26 1.86 9.14 1.86 9.14 3.58 11.02 3.58
                 11.02 2.64 13.10 2.64 ;
        POLYGON  12.24 1.54 10.06 1.54 10.06 2.54 10.60 2.54 10.60 2.86
                 9.74 2.86 9.74 1.22 12.24 1.22 ;
        POLYGON  7.86 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 7.86 4.22 ;
        RECT  6.66 1.22 7.66 1.54 ;
        RECT  5.54 3.58 6.54 3.90 ;
        RECT  5.28 1.22 6.28 1.54 ;
        POLYGON  5.08 3.90 4.62 3.90 4.62 2.40 3.68 2.40 3.68 3.08 2.14 3.08
                 2.14 3.90 1.82 3.90 1.82 3.08 0.80 3.08 0.80 2.72 1.12 2.72
                 1.12 2.76 3.36 2.76 3.36 2.08 4.58 2.08 4.58 1.22 4.90 1.22
                 4.90 2.08 4.94 2.08 4.94 3.58 5.08 3.58 ;
        POLYGON  4.30 3.90 2.50 3.90 2.50 3.58 3.98 3.58 3.98 3.36 4.30 3.36 ;
        RECT  3.20 1.22 4.20 1.54 ;
        RECT  1.58 1.22 2.82 1.54 ;
    END
END dffprqb_2

MACRO dffprqb_1
    CLASS CORE ;
    FOREIGN dffprqb_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 20.48 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  7.84 2.72 8.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.08 3.04 2.44 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.58  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.32 4.54 19.92 4.54 19.92 4.22 20.00 4.22 20.00 1.54
                 19.92 1.54 19.92 1.22 20.32 1.22 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.22  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 2.08 2.44 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 0.90 19.40 0.90 19.40 1.54 19.08 1.54 19.08 0.90
                 17.78 0.90 17.78 1.54 17.46 1.54 17.46 0.90 8.36 0.90
                 8.36 1.54 8.04 1.54 8.04 0.90 1.20 0.90 1.20 1.54 0.88 1.54
                 0.88 0.90 0.00 0.90 0.00 -0.90 20.48 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 6.66 0.00 6.66 0.00 4.86 16.08 4.86 16.08 4.12
                 16.40 4.12 16.40 4.86 17.58 4.86 17.58 4.56 17.90 4.56
                 17.90 4.86 20.48 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  19.62 3.93 19.20 4.35 18.28 4.35 18.28 3.16 16.14 3.16
                 16.14 2.84 18.28 2.84 18.28 1.54 18.16 1.54 18.16 1.22
                 18.60 1.22 18.60 4.03 19.06 4.03 19.30 3.79 19.30 2.46
                 19.26 2.46 19.26 2.14 19.62 2.14 ;
        POLYGON  17.96 2.52 15.82 2.52 15.82 3.48 17.08 3.48 17.08 4.54
                 16.76 4.54 16.76 3.80 14.46 3.80 14.22 4.04 14.22 4.54
                 13.90 4.54 13.90 3.90 14.32 3.48 15.50 3.48 15.50 2.52
                 14.76 2.52 14.00 1.76 14.00 1.22 14.32 1.22 14.32 1.62
                 14.90 2.20 17.96 2.20 ;
        RECT  16.08 1.22 17.08 1.54 ;
        RECT  14.70 1.22 15.70 1.54 ;
        RECT  14.60 4.12 15.70 4.44 ;
        POLYGON  14.06 2.60 13.74 2.60 13.74 3.24 13.08 3.90 11.98 3.90
                 11.98 4.54 8.18 4.54 8.18 4.05 8.03 3.90 6.86 3.90 6.86 3.26
                 5.90 3.26 5.90 2.94 7.18 2.94 7.18 3.58 8.17 3.58 8.50 3.91
                 8.50 4.22 11.66 4.22 11.66 3.58 12.94 3.58 13.42 3.10
                 13.42 2.50 13.10 2.18 10.38 2.18 10.38 1.86 13.24 1.86
                 13.66 2.28 14.06 2.28 ;
        RECT  12.62 1.22 13.62 1.54 ;
        RECT  12.52 4.22 13.52 4.54 ;
        POLYGON  13.10 2.96 11.34 2.96 11.34 3.90 8.82 3.90 8.82 2.18 5.58 2.18
                 5.58 3.26 5.26 3.26 5.26 1.86 9.14 1.86 9.14 3.58 11.02 3.58
                 11.02 2.64 13.10 2.64 ;
        POLYGON  12.24 1.54 10.06 1.54 10.06 2.54 10.60 2.54 10.60 2.86
                 9.74 2.86 9.74 1.22 12.24 1.22 ;
        POLYGON  7.86 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 7.86 4.22 ;
        RECT  6.66 1.22 7.66 1.54 ;
        RECT  5.54 3.58 6.54 3.90 ;
        RECT  5.28 1.22 6.28 1.54 ;
        POLYGON  5.08 3.90 4.62 3.90 4.62 2.40 3.68 2.40 3.68 3.08 2.14 3.08
                 2.14 3.90 1.82 3.90 1.82 3.08 0.80 3.08 0.80 2.72 1.12 2.72
                 1.12 2.76 3.36 2.76 3.36 2.08 4.58 2.08 4.58 1.22 4.90 1.22
                 4.90 2.08 4.94 2.08 4.94 3.58 5.08 3.58 ;
        POLYGON  4.30 3.90 2.50 3.90 2.50 3.58 3.98 3.58 3.98 3.36 4.30 3.36 ;
        RECT  3.20 1.22 4.20 1.54 ;
        RECT  1.58 1.22 2.82 1.54 ;
    END
END dffprqb_1

MACRO dffprq_4
    CLASS CORE ;
    FOREIGN dffprq_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  7.84 2.72 8.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.08 3.04 2.44 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.96 3.04 20.80 3.04 20.80 4.54 20.48 4.54 20.48 3.04
                 19.40 3.04 19.40 4.54 19.08 4.54 19.08 1.22 19.40 1.22
                 19.40 2.72 20.48 2.72 20.48 1.22 20.80 1.22 20.80 2.72
                 20.96 2.72 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.30  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 2.08 2.44 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 0.90 20.10 0.90 20.10 1.54 19.78 1.54 19.78 0.90
                 17.78 0.90 17.78 1.54 17.46 1.54 17.46 0.90 8.36 0.90
                 8.36 1.54 8.04 1.54 8.04 0.90 1.20 0.90 1.20 1.54 0.88 1.54
                 0.88 0.90 0.00 0.90 0.00 -0.90 21.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 6.66 0.00 6.66 0.00 4.86 16.08 4.86 16.08 4.12
                 16.40 4.12 16.40 4.86 17.58 4.86 17.58 4.56 17.90 4.56
                 17.90 4.86 19.78 4.86 19.78 3.58 20.10 3.58 20.10 4.86
                 21.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  18.72 4.54 18.28 4.54 18.28 3.16 16.14 3.16 16.14 2.84
                 18.28 2.84 18.28 1.54 18.16 1.54 18.16 1.22 18.60 1.22
                 18.60 4.22 18.72 4.22 ;
        POLYGON  17.96 2.52 15.82 2.52 15.82 3.48 17.08 3.48 17.08 4.54
                 16.76 4.54 16.76 3.80 14.46 3.80 14.22 4.04 14.22 4.54
                 13.90 4.54 13.90 3.90 14.32 3.48 15.50 3.48 15.50 2.52
                 14.76 2.52 14.00 1.76 14.00 1.22 14.32 1.22 14.32 1.62
                 14.90 2.20 17.96 2.20 ;
        RECT  16.08 1.22 17.08 1.54 ;
        RECT  14.70 1.22 15.70 1.54 ;
        RECT  14.60 4.12 15.70 4.44 ;
        RECT  12.62 1.22 13.62 1.54 ;
        RECT  12.52 4.22 13.52 4.54 ;
        POLYGON  13.10 2.96 11.34 2.96 11.34 3.90 8.82 3.90 8.82 2.18 5.58 2.18
                 5.58 3.26 5.26 3.26 5.26 1.86 9.14 1.86 9.14 3.58 11.02 3.58
                 11.02 2.64 13.10 2.64 ;
        POLYGON  12.24 1.54 10.06 1.54 10.06 2.54 10.60 2.54 10.60 2.86
                 9.74 2.86 9.74 1.22 12.24 1.22 ;
        POLYGON  7.86 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 7.86 4.22 ;
        RECT  6.66 1.22 7.66 1.54 ;
        RECT  5.54 3.58 6.54 3.90 ;
        RECT  5.28 1.22 6.28 1.54 ;
        POLYGON  5.08 3.90 4.62 3.90 4.62 2.40 3.68 2.40 3.68 3.08 2.14 3.08
                 2.14 3.90 1.82 3.90 1.82 3.08 0.80 3.08 0.80 2.72 1.12 2.72
                 1.12 2.76 3.36 2.76 3.36 2.08 4.58 2.08 4.58 1.22 4.90 1.22
                 4.90 2.08 4.94 2.08 4.94 3.58 5.08 3.58 ;
        POLYGON  4.30 3.90 2.50 3.90 2.50 3.58 3.98 3.58 3.98 3.36 4.30 3.36 ;
        RECT  3.20 1.22 4.20 1.54 ;
        RECT  1.58 1.22 2.82 1.54 ;
        POLYGON  14.06 2.60 13.74 2.60 13.74 3.24 13.08 3.90 11.98 3.90
                 11.98 4.54 8.18 4.54 8.18 4.05 8.03 3.90 6.86 3.90 6.86 3.26
                 5.90 3.26 5.90 2.94 7.18 2.94 7.18 3.58 8.17 3.58 8.50 3.91
                 8.50 4.22 11.66 4.22 11.66 3.58 12.94 3.58 13.42 3.10
                 13.42 2.50 13.10 2.18 10.38 2.18 10.38 1.86 13.24 1.86
                 13.66 2.28 14.06 2.28 ;
    END
END dffprq_4

MACRO dffprq_2
    CLASS CORE ;
    FOREIGN dffprq_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 20.48 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  7.84 2.72 8.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.08 3.04 2.44 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.32 3.04 20.10 3.04 20.10 4.54 19.78 4.54 19.78 1.64
                 20.10 1.64 20.10 2.72 20.32 2.72 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.22  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 2.08 2.44 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 0.90 19.40 0.90 19.40 1.96 19.08 1.96 19.08 0.90
                 17.78 0.90 17.78 1.54 17.46 1.54 17.46 0.90 8.36 0.90
                 8.36 1.54 8.04 1.54 8.04 0.90 1.20 0.90 1.20 1.54 0.88 1.54
                 0.88 0.90 0.00 0.90 0.00 -0.90 20.48 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 6.66 0.00 6.66 0.00 4.86 16.08 4.86 16.08 4.12
                 16.40 4.12 16.40 4.86 17.58 4.86 17.58 4.56 17.90 4.56
                 17.90 4.86 19.08 4.86 19.08 4.22 19.40 4.22 19.40 4.86
                 20.48 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  18.72 4.54 18.28 4.54 18.28 3.16 16.14 3.16 16.14 2.84
                 18.28 2.84 18.28 1.54 18.16 1.54 18.16 1.22 18.60 1.22
                 18.60 4.22 18.72 4.22 ;
        POLYGON  17.96 2.52 15.82 2.52 15.82 3.48 17.08 3.48 17.08 4.54
                 16.76 4.54 16.76 3.80 14.46 3.80 14.22 4.04 14.22 4.54
                 13.90 4.54 13.90 3.90 14.32 3.48 15.50 3.48 15.50 2.52
                 14.76 2.52 14.00 1.76 14.00 1.22 14.32 1.22 14.32 1.62
                 14.90 2.20 17.96 2.20 ;
        RECT  16.08 1.22 17.08 1.54 ;
        RECT  14.70 1.22 15.70 1.54 ;
        RECT  14.60 4.12 15.70 4.44 ;
        POLYGON  14.06 2.60 13.74 2.60 13.74 3.24 13.08 3.90 11.98 3.90
                 11.98 4.54 8.18 4.54 8.18 4.05 8.03 3.90 6.86 3.90 6.86 3.26
                 5.90 3.26 5.90 2.94 7.18 2.94 7.18 3.58 8.17 3.58 8.50 3.91
                 8.50 4.22 11.66 4.22 11.66 3.58 12.94 3.58 13.42 3.10
                 13.42 2.50 13.10 2.18 10.38 2.18 10.38 1.86 13.24 1.86
                 13.66 2.28 14.06 2.28 ;
        RECT  12.62 1.22 13.62 1.54 ;
        RECT  12.52 4.22 13.52 4.54 ;
        POLYGON  13.10 2.96 11.34 2.96 11.34 3.90 8.82 3.90 8.82 2.18 5.58 2.18
                 5.58 3.26 5.26 3.26 5.26 1.86 9.14 1.86 9.14 3.58 11.02 3.58
                 11.02 2.64 13.10 2.64 ;
        POLYGON  12.24 1.54 10.06 1.54 10.06 2.54 10.60 2.54 10.60 2.86
                 9.74 2.86 9.74 1.22 12.24 1.22 ;
        POLYGON  7.86 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 7.86 4.22 ;
        RECT  6.66 1.22 7.66 1.54 ;
        RECT  5.54 3.58 6.54 3.90 ;
        RECT  5.28 1.22 6.28 1.54 ;
        POLYGON  5.08 3.90 4.62 3.90 4.62 2.40 3.68 2.40 3.68 3.08 2.14 3.08
                 2.14 3.90 1.82 3.90 1.82 3.08 0.80 3.08 0.80 2.72 1.12 2.72
                 1.12 2.76 3.36 2.76 3.36 2.08 4.58 2.08 4.58 1.22 4.90 1.22
                 4.90 2.08 4.94 2.08 4.94 3.58 5.08 3.58 ;
        POLYGON  4.30 3.90 2.50 3.90 2.50 3.58 3.98 3.58 3.98 3.36 4.30 3.36 ;
        RECT  3.20 1.22 4.20 1.54 ;
        RECT  1.58 1.22 2.82 1.54 ;
    END
END dffprq_2

MACRO dffprq_1
    CLASS CORE ;
    FOREIGN dffprq_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 20.48 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  7.84 2.72 8.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.08 3.04 2.44 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.32 3.04 20.10 3.04 20.10 4.30 19.78 4.30 19.78 1.22
                 20.10 1.22 20.10 2.72 20.32 2.72 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.22  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 2.08 2.44 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 0.90 19.40 0.90 19.40 1.54 19.08 1.54 19.08 0.90
                 17.78 0.90 17.78 1.54 17.46 1.54 17.46 0.90 8.36 0.90
                 8.36 1.54 8.04 1.54 8.04 0.90 1.20 0.90 1.20 1.54 0.88 1.54
                 0.88 0.90 0.00 0.90 0.00 -0.90 20.48 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 6.66 0.00 6.66 0.00 4.86 16.08 4.86 16.08 4.12
                 16.40 4.12 16.40 4.86 17.58 4.86 17.58 4.56 17.90 4.56
                 17.90 4.86 19.08 4.86 19.08 4.06 19.40 4.06 19.40 4.86
                 20.48 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  18.72 4.54 18.28 4.54 18.28 3.16 16.14 3.16 16.14 2.84
                 18.28 2.84 18.28 1.54 18.16 1.54 18.16 1.22 18.60 1.22
                 18.60 4.22 18.72 4.22 ;
        POLYGON  17.96 2.52 15.82 2.52 15.82 3.48 17.08 3.48 17.08 4.54
                 16.76 4.54 16.76 3.80 14.46 3.80 14.22 4.04 14.22 4.54
                 13.90 4.54 13.90 3.90 14.32 3.48 15.50 3.48 15.50 2.52
                 14.76 2.52 14.00 1.76 14.00 1.22 14.32 1.22 14.32 1.62
                 14.90 2.20 17.96 2.20 ;
        RECT  16.08 1.22 17.08 1.54 ;
        RECT  14.70 1.22 15.70 1.54 ;
        RECT  14.60 4.12 15.70 4.44 ;
        POLYGON  14.06 2.60 13.74 2.60 13.74 3.24 13.08 3.90 11.98 3.90
                 11.98 4.54 8.18 4.54 8.18 4.05 8.03 3.90 6.86 3.90 6.86 3.26
                 5.90 3.26 5.90 2.94 7.18 2.94 7.18 3.58 8.17 3.58 8.50 3.91
                 8.50 4.22 11.66 4.22 11.66 3.58 12.94 3.58 13.42 3.10
                 13.42 2.50 13.10 2.18 10.38 2.18 10.38 1.86 13.24 1.86
                 13.66 2.28 14.06 2.28 ;
        RECT  12.62 1.22 13.62 1.54 ;
        RECT  12.52 4.22 13.52 4.54 ;
        POLYGON  13.10 2.96 11.34 2.96 11.34 3.90 8.82 3.90 8.82 2.18 5.58 2.18
                 5.58 3.26 5.26 3.26 5.26 1.86 9.14 1.86 9.14 3.58 11.02 3.58
                 11.02 2.64 13.10 2.64 ;
        POLYGON  12.24 1.54 10.06 1.54 10.06 2.54 10.60 2.54 10.60 2.86
                 9.74 2.86 9.74 1.22 12.24 1.22 ;
        POLYGON  7.86 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 7.86 4.22 ;
        RECT  6.66 1.22 7.66 1.54 ;
        RECT  5.54 3.58 6.54 3.90 ;
        RECT  5.28 1.22 6.28 1.54 ;
        POLYGON  5.08 3.90 4.62 3.90 4.62 2.40 3.68 2.40 3.68 3.08 2.14 3.08
                 2.14 3.90 1.82 3.90 1.82 3.08 0.80 3.08 0.80 2.72 1.12 2.72
                 1.12 2.76 3.36 2.76 3.36 2.08 4.58 2.08 4.58 1.22 4.90 1.22
                 4.90 2.08 4.94 2.08 4.94 3.58 5.08 3.58 ;
        POLYGON  4.30 3.90 2.50 3.90 2.50 3.58 3.98 3.58 3.98 3.36 4.30 3.36 ;
        RECT  3.20 1.22 4.20 1.54 ;
        RECT  1.58 1.22 2.82 1.54 ;
    END
END dffprq_1

MACRO dffpr_4
    CLASS CORE ;
    FOREIGN dffpr_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  7.84 2.72 8.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.08 3.04 2.44 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  21.05 3.25 19.32 3.25 19.32 2.93 20.64 2.93 20.64 1.54
                 18.84 1.54 18.84 1.22 20.96 1.22 20.96 2.71 21.05 2.71 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  23.52 4.53 21.41 4.53 21.41 4.21 23.20 4.21 23.20 1.90
                 21.41 1.90 21.41 1.58 23.52 1.58 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.22  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 2.08 2.44 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  23.68 0.90 22.43 0.90 22.43 1.23 22.11 1.23 22.11 0.90
                 17.78 0.90 17.78 1.54 17.46 1.54 17.46 0.90 8.36 0.90
                 8.36 1.54 8.04 1.54 8.04 0.90 1.20 0.90 1.20 1.54 0.88 1.54
                 0.88 0.90 0.00 0.90 0.00 -0.90 23.68 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  23.68 6.66 0.00 6.66 0.00 4.86 16.08 4.86 16.08 4.20
                 16.40 4.20 16.40 4.86 17.58 4.86 17.58 4.56 17.90 4.56
                 17.90 4.86 19.99 4.86 19.99 4.81 20.37 4.81 20.37 4.86
                 23.68 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  22.43 3.89 18.72 3.89 18.72 4.54 18.40 4.54 18.40 3.22
                 16.14 3.22 16.14 2.90 18.28 2.90 18.28 2.02 18.16 2.02
                 18.16 1.22 18.48 1.22 18.48 1.76 18.60 1.76 18.60 2.90
                 18.72 2.90 18.72 3.57 22.11 3.57 22.11 2.65 22.07 2.65
                 22.07 2.33 22.43 2.33 ;
        POLYGON  17.94 2.58 15.82 2.58 15.82 3.54 17.08 3.54 17.08 4.54
                 16.76 4.54 16.76 3.86 14.40 3.86 14.22 4.04 14.22 4.54
                 13.90 4.54 13.90 3.90 14.26 3.54 15.50 3.54 15.50 2.58
                 14.82 2.58 14.00 1.76 14.00 1.22 14.32 1.22 14.32 1.62
                 14.96 2.26 17.94 2.26 ;
        RECT  16.08 1.22 17.08 1.54 ;
        RECT  14.70 1.22 15.70 1.54 ;
        RECT  14.60 4.20 15.70 4.52 ;
        POLYGON  14.06 2.60 13.74 2.60 13.74 3.24 13.08 3.90 11.98 3.90
                 11.98 4.54 8.18 4.54 8.18 4.05 8.03 3.90 6.86 3.90 6.86 3.26
                 5.90 3.26 5.90 2.94 7.18 2.94 7.18 3.58 8.17 3.58 8.50 3.91
                 8.50 4.22 11.66 4.22 11.66 3.58 12.94 3.58 13.42 3.10
                 13.42 2.50 13.10 2.18 10.38 2.18 10.38 1.86 13.24 1.86
                 13.66 2.28 14.06 2.28 ;
        RECT  12.62 1.22 13.62 1.54 ;
        RECT  12.52 4.22 13.52 4.54 ;
        POLYGON  13.10 2.96 11.34 2.96 11.34 3.90 8.82 3.90 8.82 2.18 5.58 2.18
                 5.58 3.26 5.26 3.26 5.26 1.86 9.14 1.86 9.14 3.58 11.02 3.58
                 11.02 2.64 13.10 2.64 ;
        POLYGON  12.24 1.54 10.06 1.54 10.06 2.54 10.60 2.54 10.60 2.86
                 9.74 2.86 9.74 1.22 12.24 1.22 ;
        POLYGON  7.86 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 7.86 4.22 ;
        RECT  6.66 1.22 7.66 1.54 ;
        RECT  5.54 3.58 6.54 3.90 ;
        RECT  5.28 1.22 6.28 1.54 ;
        POLYGON  5.08 3.90 4.62 3.90 4.62 2.40 3.68 2.40 3.68 3.08 2.14 3.08
                 2.14 3.90 1.82 3.90 1.82 3.08 0.80 3.08 0.80 2.72 1.12 2.72
                 1.12 2.76 3.36 2.76 3.36 2.08 4.58 2.08 4.58 1.22 4.90 1.22
                 4.90 2.08 4.94 2.08 4.94 3.58 5.08 3.58 ;
        POLYGON  4.30 3.90 2.50 3.90 2.50 3.58 3.98 3.58 3.98 3.36 4.30 3.36 ;
        RECT  3.20 1.22 4.20 1.54 ;
        RECT  1.58 1.22 2.82 1.54 ;
    END
END dffpr_4

MACRO dffpr_2
    CLASS CORE ;
    FOREIGN dffpr_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  7.84 2.72 8.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.08 3.04 2.44 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  19.68 3.04 19.40 3.04 19.40 3.47 19.04 3.47 19.04 1.26
                 19.40 1.26 19.40 1.58 19.36 1.58 19.36 2.72 19.68 2.72 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.19  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.96 4.54 20.62 4.54 20.62 4.22 20.64 4.22 20.64 1.58
                 20.62 1.58 20.62 1.26 20.96 1.26 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.22  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 2.08 2.44 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 0.90 20.10 0.90 20.10 1.58 19.78 1.58 19.78 0.90
                 17.78 0.90 17.78 1.54 17.46 1.54 17.46 0.90 8.36 0.90
                 8.36 1.54 8.04 1.54 8.04 0.90 1.20 0.90 1.20 1.54 0.88 1.54
                 0.88 0.90 0.00 0.90 0.00 -0.90 21.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 6.66 0.00 6.66 0.00 4.86 16.08 4.86 16.08 4.12
                 16.40 4.12 16.40 4.86 17.58 4.86 17.58 4.56 17.90 4.56
                 17.90 4.86 21.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.32 3.91 19.69 4.54 18.28 4.54 18.28 3.16 16.14 3.16
                 16.14 2.84 18.28 2.84 18.28 1.54 18.16 1.54 18.16 1.22
                 18.60 1.22 18.60 4.22 19.54 4.22 20.00 3.76 20.00 2.46
                 19.96 2.46 19.96 2.14 20.32 2.14 ;
        POLYGON  17.96 2.52 15.82 2.52 15.82 3.48 17.08 3.48 17.08 4.54
                 16.76 4.54 16.76 3.80 14.46 3.80 14.22 4.04 14.22 4.54
                 13.90 4.54 13.90 3.90 14.32 3.48 15.50 3.48 15.50 2.52
                 14.76 2.52 14.00 1.76 14.00 1.22 14.32 1.22 14.32 1.62
                 14.90 2.20 17.96 2.20 ;
        RECT  16.08 1.22 17.08 1.54 ;
        RECT  14.70 1.22 15.70 1.54 ;
        RECT  14.60 4.12 15.70 4.44 ;
        POLYGON  14.06 2.60 13.74 2.60 13.74 3.24 13.08 3.90 11.98 3.90
                 11.98 4.54 8.18 4.54 8.18 4.05 8.03 3.90 6.86 3.90 6.86 3.26
                 5.90 3.26 5.90 2.94 7.18 2.94 7.18 3.58 8.17 3.58 8.50 3.91
                 8.50 4.22 11.66 4.22 11.66 3.58 12.94 3.58 13.42 3.10
                 13.42 2.50 13.10 2.18 10.38 2.18 10.38 1.86 13.24 1.86
                 13.66 2.28 14.06 2.28 ;
        RECT  12.62 1.22 13.62 1.54 ;
        RECT  12.52 4.22 13.52 4.54 ;
        POLYGON  13.10 2.96 11.34 2.96 11.34 3.90 8.82 3.90 8.82 2.18 5.58 2.18
                 5.58 3.26 5.26 3.26 5.26 1.86 9.14 1.86 9.14 3.58 11.02 3.58
                 11.02 2.64 13.10 2.64 ;
        POLYGON  12.24 1.54 10.06 1.54 10.06 2.54 10.60 2.54 10.60 2.86
                 9.74 2.86 9.74 1.22 12.24 1.22 ;
        POLYGON  7.86 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 7.86 4.22 ;
        RECT  6.66 1.22 7.66 1.54 ;
        RECT  5.54 3.58 6.54 3.90 ;
        RECT  5.28 1.22 6.28 1.54 ;
        POLYGON  5.08 3.90 4.62 3.90 4.62 2.40 3.68 2.40 3.68 3.08 2.14 3.08
                 2.14 3.90 1.82 3.90 1.82 3.08 0.80 3.08 0.80 2.72 1.12 2.72
                 1.12 2.76 3.36 2.76 3.36 2.08 4.58 2.08 4.58 1.22 4.90 1.22
                 4.90 2.08 4.94 2.08 4.94 3.58 5.08 3.58 ;
        POLYGON  4.30 3.90 2.50 3.90 2.50 3.58 3.98 3.58 3.98 3.36 4.30 3.36 ;
        RECT  3.20 1.22 4.20 1.54 ;
        RECT  1.58 1.22 2.82 1.54 ;
    END
END dffpr_2

MACRO dffpr_1
    CLASS CORE ;
    FOREIGN dffpr_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  7.84 2.72 8.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.08 3.04 2.44 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.21  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  19.68 3.04 19.36 3.04 19.36 3.58 19.40 3.58 19.40 3.90
                 19.04 3.90 19.04 1.22 19.40 1.22 19.40 1.54 19.36 1.54
                 19.36 2.72 19.68 2.72 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.96 4.54 20.62 4.54 20.62 4.22 20.64 4.22 20.64 1.54
                 20.62 1.54 20.62 1.22 20.96 1.22 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.22  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 2.08 2.44 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 0.90 20.10 0.90 20.10 1.54 19.78 1.54 19.78 0.90
                 17.78 0.90 17.78 1.54 17.46 1.54 17.46 0.90 8.36 0.90
                 8.36 1.54 8.04 1.54 8.04 0.90 1.20 0.90 1.20 1.54 0.88 1.54
                 0.88 0.90 0.00 0.90 0.00 -0.90 21.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 6.66 0.00 6.66 0.00 4.86 16.08 4.86 16.08 4.12
                 16.40 4.12 16.40 4.86 17.58 4.86 17.58 4.56 17.90 4.56
                 17.90 4.86 21.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.32 3.91 19.69 4.54 18.28 4.54 18.28 3.16 16.14 3.16
                 16.14 2.84 18.28 2.84 18.28 1.54 18.16 1.54 18.16 1.22
                 18.60 1.22 18.60 4.22 19.54 4.22 20.00 3.76 20.00 2.46
                 19.96 2.46 19.96 2.14 20.32 2.14 ;
        POLYGON  17.96 2.52 15.82 2.52 15.82 3.48 17.08 3.48 17.08 4.54
                 16.76 4.54 16.76 3.80 14.46 3.80 14.22 4.04 14.22 4.54
                 13.90 4.54 13.90 3.90 14.32 3.48 15.50 3.48 15.50 2.52
                 14.76 2.52 14.00 1.76 14.00 1.22 14.32 1.22 14.32 1.62
                 14.90 2.20 17.96 2.20 ;
        RECT  16.08 1.22 17.08 1.54 ;
        RECT  14.70 1.22 15.70 1.54 ;
        RECT  14.60 4.12 15.70 4.44 ;
        POLYGON  14.06 2.60 13.74 2.60 13.74 3.24 13.08 3.90 11.98 3.90
                 11.98 4.54 8.18 4.54 8.18 4.05 8.03 3.90 6.86 3.90 6.86 3.26
                 5.90 3.26 5.90 2.94 7.18 2.94 7.18 3.58 8.17 3.58 8.50 3.91
                 8.50 4.22 11.66 4.22 11.66 3.58 12.94 3.58 13.42 3.10
                 13.42 2.50 13.10 2.18 10.38 2.18 10.38 1.86 13.24 1.86
                 13.66 2.28 14.06 2.28 ;
        RECT  12.62 1.22 13.62 1.54 ;
        RECT  12.52 4.22 13.52 4.54 ;
        POLYGON  13.10 2.96 11.34 2.96 11.34 3.90 8.82 3.90 8.82 2.18 5.58 2.18
                 5.58 3.26 5.26 3.26 5.26 1.86 9.14 1.86 9.14 3.58 11.02 3.58
                 11.02 2.64 13.10 2.64 ;
        POLYGON  12.24 1.54 10.06 1.54 10.06 2.54 10.60 2.54 10.60 2.86
                 9.74 2.86 9.74 1.22 12.24 1.22 ;
        POLYGON  7.86 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 7.86 4.22 ;
        RECT  6.66 1.22 7.66 1.54 ;
        RECT  5.54 3.58 6.54 3.90 ;
        RECT  5.28 1.22 6.28 1.54 ;
        POLYGON  5.08 3.90 4.62 3.90 4.62 2.40 3.68 2.40 3.68 3.08 2.14 3.08
                 2.14 3.90 1.82 3.90 1.82 3.08 0.80 3.08 0.80 2.72 1.12 2.72
                 1.12 2.76 3.36 2.76 3.36 2.08 4.58 2.08 4.58 1.22 4.90 1.22
                 4.90 2.08 4.94 2.08 4.94 3.58 5.08 3.58 ;
        POLYGON  4.30 3.90 2.50 3.90 2.50 3.58 3.98 3.58 3.98 3.36 4.30 3.36 ;
        RECT  3.20 1.22 4.20 1.54 ;
        RECT  1.58 1.22 2.82 1.54 ;
    END
END dffpr_1

MACRO dffpqb_4
    CLASS CORE ;
    FOREIGN dffpqb_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.64 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.03 3.46 8.84 3.46 8.80 3.50 8.80 3.90 8.48 3.90 8.48 3.36
                 8.70 3.14 9.03 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.42 2.08 2.06 2.40 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.48 4.53 14.49 4.53 14.49 4.21 16.16 4.21 16.16 1.90
                 14.49 1.90 14.49 1.58 16.48 1.58 ;
        END
    END qb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 0.90 15.52 0.90 15.52 1.24 15.18 1.24 15.18 0.90
                 13.14 0.90 13.14 1.54 12.82 1.54 12.82 0.90 6.07 0.90
                 6.07 1.14 5.75 1.14 5.75 0.90 1.32 0.90 1.32 1.34 1.00 1.34
                 1.00 0.90 0.00 0.90 0.00 -0.90 16.64 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 6.66 0.00 6.66 0.00 4.86 5.94 4.86 5.94 3.74 6.26 3.74
                 6.26 4.86 12.93 4.86 12.93 3.96 13.25 3.96 13.25 4.86
                 16.64 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  15.51 3.89 13.64 3.89 13.64 3.53 13.57 3.53 13.57 3.18
                 12.42 3.18 12.42 2.86 13.57 2.86 13.57 1.22 13.89 1.22
                 13.89 3.21 13.96 3.21 13.96 3.57 15.19 3.57 15.19 2.34
                 15.51 2.34 ;
        POLYGON  13.25 2.47 12.93 2.47 12.93 2.28 11.03 2.28 11.03 4.54
                 10.71 4.54 10.71 2.28 10.27 1.84 10.27 1.22 10.59 1.22
                 10.59 1.70 10.85 1.96 13.25 1.96 ;
        RECT  11.49 3.96 12.49 4.28 ;
        RECT  11.09 1.22 12.39 1.54 ;
        POLYGON  10.39 3.90 9.33 3.90 9.33 3.58 10.07 3.58 10.07 2.60 9.65 2.18
                 7.51 2.18 7.29 2.40 7.29 2.58 6.97 2.58 6.97 2.26 7.37 1.86
                 9.79 1.86 10.39 2.46 ;
        RECT  7.37 4.22 10.33 4.54 ;
        RECT  7.13 1.22 9.77 1.54 ;
        POLYGON  9.51 2.82 8.55 2.82 7.95 3.42 7.09 3.42 7.09 3.90 6.77 3.90
                 6.77 3.42 6.33 3.42 6.33 2.32 3.88 2.32 3.88 2.00 6.33 2.00
                 6.33 1.66 6.45 1.66 6.45 1.22 6.77 1.22 6.77 1.99 6.65 1.99
                 6.65 3.10 7.81 3.10 8.41 2.50 9.51 2.50 ;
        RECT  4.41 3.46 5.45 3.78 ;
        RECT  4.00 1.22 5.37 1.54 ;
        POLYGON  5.09 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 5.09 4.22 ;
        POLYGON  4.03 3.90 3.30 3.90 3.30 3.04 0.80 3.04 0.80 2.66 1.12 2.66
                 1.12 2.72 2.92 2.72 2.92 2.00 3.30 1.62 3.30 1.22 3.62 1.22
                 3.62 1.76 3.24 2.14 3.24 2.72 3.62 2.72 3.62 3.58 4.03 3.58 ;
        RECT  1.82 1.22 2.92 1.54 ;
        RECT  1.82 3.58 2.92 3.90 ;
    END
END dffpqb_4

MACRO dffpqb_2
    CLASS CORE ;
    FOREIGN dffpqb_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.00 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.03 3.46 8.84 3.46 8.80 3.50 8.80 3.90 8.48 3.90 8.48 3.36
                 8.70 3.14 9.03 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.42 2.08 2.06 2.40 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  15.84 4.54 15.19 4.54 15.19 4.22 15.52 4.22 15.52 1.77
                 15.19 1.77 15.19 1.45 15.84 1.45 ;
        END
    END qb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 0.90 14.81 0.90 14.81 1.24 14.49 1.24 14.49 0.90
                 13.19 0.90 13.19 1.14 12.87 1.14 12.87 0.90 6.07 0.90
                 6.07 1.14 5.75 1.14 5.75 0.90 1.32 0.90 1.32 1.34 1.00 1.34
                 1.00 0.90 0.00 0.90 0.00 -0.90 16.00 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 6.66 0.00 6.66 0.00 4.86 5.94 4.86 5.94 3.74 6.26 3.74
                 6.26 4.86 12.93 4.86 12.93 3.96 13.25 3.96 13.25 4.86
                 16.00 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  14.99 3.84 14.74 3.84 14.74 4.54 13.57 4.54 13.57 3.18
                 12.59 3.18 12.59 2.86 13.57 2.86 13.57 1.22 13.89 1.22
                 13.89 4.22 14.42 4.22 14.42 3.52 14.67 3.52 14.67 2.14
                 14.99 2.14 ;
        POLYGON  13.25 2.47 12.93 2.47 12.93 2.28 11.03 2.28 11.03 4.54
                 10.71 4.54 10.71 2.28 10.27 1.84 10.27 1.22 10.59 1.22
                 10.59 1.70 10.85 1.96 13.25 1.96 ;
        RECT  11.49 3.96 12.49 4.28 ;
        RECT  11.09 1.22 12.39 1.54 ;
        POLYGON  10.39 3.90 9.33 3.90 9.33 3.58 10.07 3.58 10.07 2.60 9.65 2.18
                 7.51 2.18 7.29 2.40 7.29 2.58 6.97 2.58 6.97 2.26 7.37 1.86
                 9.79 1.86 10.39 2.46 ;
        RECT  7.37 4.22 10.33 4.54 ;
        RECT  7.13 1.22 9.77 1.54 ;
        POLYGON  9.51 2.82 8.55 2.82 7.95 3.42 7.09 3.42 7.09 3.90 6.77 3.90
                 6.77 3.42 6.33 3.42 6.33 2.32 3.88 2.32 3.88 2.00 6.33 2.00
                 6.33 1.66 6.45 1.66 6.45 1.22 6.77 1.22 6.77 1.99 6.65 1.99
                 6.65 3.10 7.81 3.10 8.41 2.50 9.51 2.50 ;
        RECT  4.41 3.46 5.45 3.78 ;
        RECT  4.00 1.22 5.37 1.54 ;
        POLYGON  5.09 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 5.09 4.22 ;
        POLYGON  4.03 3.90 3.30 3.90 3.30 3.04 0.80 3.04 0.80 2.66 1.12 2.66
                 1.12 2.72 2.92 2.72 2.92 2.00 3.30 1.62 3.30 1.22 3.62 1.22
                 3.62 1.76 3.24 2.14 3.24 2.72 3.62 2.72 3.62 3.58 4.03 3.58 ;
        RECT  1.82 1.22 2.92 1.54 ;
        RECT  1.82 3.58 2.92 3.90 ;
    END
END dffpqb_2

MACRO dffpqb_1
    CLASS CORE ;
    FOREIGN dffpqb_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.00 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.03 3.46 8.84 3.46 8.80 3.50 8.80 3.90 8.48 3.90 8.48 3.36
                 8.70 3.14 9.03 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.42 2.08 2.06 2.40 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  15.84 4.54 15.27 4.54 15.27 4.22 15.52 4.22 15.52 1.55
                 14.95 1.55 14.95 1.23 15.84 1.23 ;
        END
    END qb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 0.90 14.57 0.90 14.57 1.24 14.25 1.24 14.25 0.90
                 13.19 0.90 13.19 1.14 12.87 1.14 12.87 0.90 6.07 0.90
                 6.07 1.14 5.75 1.14 5.75 0.90 1.32 0.90 1.32 1.34 1.00 1.34
                 1.00 0.90 0.00 0.90 0.00 -0.90 16.00 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 6.66 0.00 6.66 0.00 4.86 5.94 4.86 5.94 3.74 6.26 3.74
                 6.26 4.86 12.93 4.86 12.93 3.96 13.25 3.96 13.25 4.86
                 16.00 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  14.75 4.54 13.57 4.54 13.57 3.18 12.59 3.18 12.59 2.86
                 13.57 2.86 13.57 1.22 13.89 1.22 13.89 4.22 14.43 4.22
                 14.43 2.46 14.41 2.46 14.41 2.14 14.75 2.14 ;
        POLYGON  13.25 2.47 12.93 2.47 12.93 2.28 11.03 2.28 11.03 4.54
                 10.71 4.54 10.71 2.28 10.27 1.84 10.27 1.22 10.59 1.22
                 10.59 1.70 10.85 1.96 13.25 1.96 ;
        RECT  11.49 3.96 12.49 4.28 ;
        RECT  11.09 1.22 12.39 1.54 ;
        POLYGON  10.39 3.90 9.33 3.90 9.33 3.58 10.07 3.58 10.07 2.60 9.65 2.18
                 7.51 2.18 7.29 2.40 7.29 2.58 6.97 2.58 6.97 2.26 7.37 1.86
                 9.79 1.86 10.39 2.46 ;
        RECT  7.37 4.22 10.33 4.54 ;
        RECT  7.13 1.22 9.77 1.54 ;
        POLYGON  9.51 2.82 8.55 2.82 7.95 3.42 7.09 3.42 7.09 3.90 6.77 3.90
                 6.77 3.42 6.33 3.42 6.33 2.32 3.88 2.32 3.88 2.00 6.33 2.00
                 6.33 1.66 6.45 1.66 6.45 1.22 6.77 1.22 6.77 1.99 6.65 1.99
                 6.65 3.10 7.81 3.10 8.41 2.50 9.51 2.50 ;
        RECT  4.41 3.46 5.45 3.78 ;
        RECT  4.00 1.22 5.37 1.54 ;
        POLYGON  5.09 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 5.09 4.22 ;
        POLYGON  4.03 3.90 3.30 3.90 3.30 3.04 0.80 3.04 0.80 2.66 1.12 2.66
                 1.12 2.72 2.92 2.72 2.92 2.00 3.30 1.62 3.30 1.22 3.62 1.22
                 3.62 1.76 3.24 2.14 3.24 2.72 3.62 2.72 3.62 3.58 4.03 3.58 ;
        RECT  1.82 1.22 2.92 1.54 ;
        RECT  1.82 3.58 2.92 3.90 ;
    END
END dffpqb_1

MACRO dffpq_4
    CLASS CORE ;
    FOREIGN dffpq_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.64 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.03 3.46 8.84 3.46 8.80 3.50 8.80 3.90 8.48 3.90 8.48 3.36
                 8.70 3.14 9.03 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.42 2.08 2.06 2.40 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.21 4.54 15.89 4.54 15.89 3.04 14.57 3.04 14.57 3.43
                 14.81 3.43 14.81 4.54 14.49 4.54 14.49 3.75 14.24 3.75
                 14.24 1.22 14.57 1.22 14.57 2.72 15.65 2.72 15.65 1.33
                 15.97 1.33 15.97 2.72 16.21 2.72 ;
        END
    END q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 0.90 15.27 0.90 15.27 1.67 14.95 1.67 14.95 0.90
                 13.19 0.90 13.19 1.14 12.87 1.14 12.87 0.90 6.07 0.90
                 6.07 1.14 5.75 1.14 5.75 0.90 1.32 0.90 1.32 1.34 1.00 1.34
                 1.00 0.90 0.00 0.90 0.00 -0.90 16.64 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 6.66 0.00 6.66 0.00 4.86 5.94 4.86 5.94 3.74 6.26 3.74
                 6.26 4.86 12.93 4.86 12.93 3.96 13.25 3.96 13.25 4.86
                 15.19 4.86 15.19 3.66 15.51 3.66 15.51 4.86 16.64 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  14.13 4.54 13.57 4.54 13.57 3.18 12.59 3.18 12.59 2.86
                 13.57 2.86 13.57 1.22 13.89 1.22 13.89 4.22 14.13 4.22 ;
        POLYGON  13.25 2.47 12.93 2.47 12.93 2.28 11.03 2.28 11.03 4.54
                 10.71 4.54 10.71 2.28 10.27 1.84 10.27 1.22 10.59 1.22
                 10.59 1.70 10.85 1.96 13.25 1.96 ;
        RECT  11.49 3.96 12.49 4.28 ;
        RECT  11.09 1.22 12.39 1.54 ;
        POLYGON  10.39 3.90 9.33 3.90 9.33 3.58 10.07 3.58 10.07 2.60 9.65 2.18
                 7.51 2.18 7.29 2.40 7.29 2.58 6.97 2.58 6.97 2.26 7.37 1.86
                 9.79 1.86 10.39 2.46 ;
        RECT  7.37 4.22 10.33 4.54 ;
        RECT  7.13 1.22 9.77 1.54 ;
        POLYGON  9.51 2.82 8.55 2.82 7.95 3.42 7.09 3.42 7.09 3.90 6.77 3.90
                 6.77 3.42 6.33 3.42 6.33 2.32 3.88 2.32 3.88 2.00 6.33 2.00
                 6.33 1.66 6.45 1.66 6.45 1.22 6.77 1.22 6.77 1.99 6.65 1.99
                 6.65 3.10 7.81 3.10 8.41 2.50 9.51 2.50 ;
        RECT  4.41 3.46 5.45 3.78 ;
        RECT  4.00 1.22 5.37 1.54 ;
        POLYGON  5.09 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 5.09 4.22 ;
        POLYGON  4.03 3.90 3.30 3.90 3.30 3.04 0.80 3.04 0.80 2.66 1.12 2.66
                 1.12 2.72 2.92 2.72 2.92 2.00 3.30 1.62 3.30 1.22 3.62 1.22
                 3.62 1.76 3.24 2.14 3.24 2.72 3.62 2.72 3.62 3.58 4.03 3.58 ;
        RECT  1.82 1.22 2.92 1.54 ;
        RECT  1.82 3.58 2.92 3.90 ;
    END
END dffpq_4

MACRO dffpq_2
    CLASS CORE ;
    FOREIGN dffpq_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.00 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.03 3.46 8.84 3.46 8.80 3.50 8.80 3.90 8.48 3.90 8.48 3.36
                 8.70 3.14 9.03 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.42 2.08 2.06 2.40 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.81 4.54 14.49 4.54 14.49 3.68 14.24 3.68 14.24 3.36
                 14.25 3.36 14.25 1.64 14.57 1.64 14.57 3.36 14.81 3.36 ;
        END
    END q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 0.90 15.27 0.90 15.27 1.24 14.95 1.24 14.95 0.90
                 13.13 0.90 13.13 1.14 12.81 1.14 12.81 0.90 6.07 0.90
                 6.07 1.14 5.75 1.14 5.75 0.90 1.32 0.90 1.32 1.34 1.00 1.34
                 1.00 0.90 0.00 0.90 0.00 -0.90 16.00 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 6.66 0.00 6.66 0.00 4.86 5.94 4.86 5.94 3.74 6.26 3.74
                 6.26 4.86 12.93 4.86 12.93 3.96 13.25 3.96 13.25 4.86
                 15.19 4.86 15.19 4.22 15.51 4.22 15.51 4.86 16.00 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  14.13 4.54 13.57 4.54 13.57 3.18 12.59 3.18 12.59 2.86
                 13.57 2.86 13.57 1.22 13.89 1.22 13.89 4.22 14.13 4.22 ;
        POLYGON  13.25 2.47 12.93 2.47 12.93 2.28 11.03 2.28 11.03 4.54
                 10.71 4.54 10.71 2.28 10.27 1.84 10.27 1.22 10.59 1.22
                 10.59 1.70 10.85 1.96 13.25 1.96 ;
        RECT  11.49 3.96 12.49 4.28 ;
        RECT  11.09 1.22 12.39 1.54 ;
        POLYGON  10.39 3.90 9.33 3.90 9.33 3.58 10.07 3.58 10.07 2.60 9.65 2.18
                 7.51 2.18 7.29 2.40 7.29 2.58 6.97 2.58 6.97 2.26 7.37 1.86
                 9.79 1.86 10.39 2.46 ;
        RECT  7.37 4.22 10.33 4.54 ;
        RECT  7.13 1.22 9.77 1.54 ;
        POLYGON  9.51 2.82 8.55 2.82 7.95 3.42 7.09 3.42 7.09 3.90 6.77 3.90
                 6.77 3.42 6.33 3.42 6.33 2.32 3.88 2.32 3.88 2.00 6.33 2.00
                 6.33 1.66 6.45 1.66 6.45 1.22 6.77 1.22 6.77 1.99 6.65 1.99
                 6.65 3.10 7.81 3.10 8.41 2.50 9.51 2.50 ;
        RECT  4.41 3.46 5.45 3.78 ;
        RECT  4.00 1.22 5.37 1.54 ;
        POLYGON  5.09 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 5.09 4.22 ;
        POLYGON  4.03 3.90 3.30 3.90 3.30 3.04 0.80 3.04 0.80 2.66 1.12 2.66
                 1.12 2.72 2.92 2.72 2.92 2.00 3.30 1.62 3.30 1.22 3.62 1.22
                 3.62 1.76 3.24 2.14 3.24 2.72 3.62 2.72 3.62 3.58 4.03 3.58 ;
        RECT  1.82 1.22 2.92 1.54 ;
        RECT  1.82 3.58 2.92 3.90 ;
    END
END dffpq_2

MACRO dffpq_1
    CLASS CORE ;
    FOREIGN dffpq_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.00 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.03 3.46 8.84 3.46 8.80 3.50 8.80 3.90 8.48 3.90 8.48 3.36
                 8.70 3.14 9.03 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.42 2.08 2.06 2.40 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.81 4.08 14.49 4.08 14.49 3.68 14.24 3.68 14.24 3.36
                 14.25 3.36 14.25 1.22 14.57 1.22 14.57 3.36 14.81 3.36 ;
        END
    END q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 0.90 15.27 0.90 15.27 1.14 14.95 1.14 14.95 0.90
                 13.13 0.90 13.13 1.14 12.81 1.14 12.81 0.90 6.07 0.90
                 6.07 1.14 5.75 1.14 5.75 0.90 1.32 0.90 1.32 1.34 1.00 1.34
                 1.00 0.90 0.00 0.90 0.00 -0.90 16.00 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 6.66 0.00 6.66 0.00 4.86 5.94 4.86 5.94 3.74 6.26 3.74
                 6.26 4.86 12.93 4.86 12.93 3.96 13.25 3.96 13.25 4.86
                 15.19 4.86 15.19 4.28 15.51 4.28 15.51 4.86 16.00 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  14.13 4.32 13.57 4.32 13.57 3.18 12.59 3.18 12.59 2.86
                 13.57 2.86 13.57 1.22 13.89 1.22 13.89 4.00 14.13 4.00 ;
        POLYGON  13.25 2.47 12.93 2.47 12.93 2.28 11.03 2.28 11.03 4.54
                 10.71 4.54 10.71 2.28 10.27 1.84 10.27 1.22 10.59 1.22
                 10.59 1.70 10.85 1.96 13.25 1.96 ;
        RECT  11.49 3.96 12.49 4.28 ;
        RECT  11.09 1.22 12.39 1.54 ;
        POLYGON  10.39 3.90 9.33 3.90 9.33 3.58 10.07 3.58 10.07 2.60 9.65 2.18
                 7.51 2.18 7.29 2.40 7.29 2.58 6.97 2.58 6.97 2.26 7.37 1.86
                 9.79 1.86 10.39 2.46 ;
        RECT  7.37 4.22 10.33 4.54 ;
        RECT  7.13 1.22 9.77 1.54 ;
        POLYGON  9.51 2.82 8.55 2.82 7.95 3.42 7.09 3.42 7.09 3.90 6.77 3.90
                 6.77 3.42 6.33 3.42 6.33 2.32 3.88 2.32 3.88 2.00 6.33 2.00
                 6.33 1.66 6.45 1.66 6.45 1.22 6.77 1.22 6.77 1.99 6.65 1.99
                 6.65 3.10 7.81 3.10 8.41 2.50 9.51 2.50 ;
        RECT  4.41 3.46 5.45 3.78 ;
        RECT  4.00 1.22 5.37 1.54 ;
        POLYGON  5.09 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 5.09 4.22 ;
        POLYGON  4.03 3.90 3.30 3.90 3.30 3.04 0.80 3.04 0.80 2.66 1.12 2.66
                 1.12 2.72 2.92 2.72 2.92 2.00 3.30 1.62 3.30 1.22 3.62 1.22
                 3.62 1.76 3.24 2.14 3.24 2.72 3.62 2.72 3.62 3.58 4.03 3.58 ;
        RECT  1.82 1.22 2.92 1.54 ;
        RECT  1.82 3.58 2.92 3.90 ;
    END
END dffpq_1

MACRO dffp_4
    CLASS CORE ;
    FOREIGN dffp_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.20 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.03 3.46 8.84 3.46 8.80 3.50 8.80 3.90 8.48 3.90 8.48 3.36
                 8.70 3.14 9.03 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.42 2.08 2.06 2.40 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.48 3.25 14.73 3.25 14.73 2.93 16.16 2.93 16.16 1.54
                 14.25 1.54 14.25 1.22 16.48 1.22 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  19.04 4.53 16.82 4.53 16.82 4.21 18.72 4.21 18.72 1.90
                 16.82 1.90 16.82 1.58 19.04 1.58 ;
        END
    END qb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  19.20 0.90 17.85 0.90 17.85 1.24 17.51 1.24 17.51 0.90
                 13.14 0.90 13.14 1.54 12.82 1.54 12.82 0.90 6.07 0.90
                 6.07 1.14 5.75 1.14 5.75 0.90 1.32 0.90 1.32 1.34 1.00 1.34
                 1.00 0.90 0.00 0.90 0.00 -0.90 19.20 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  19.20 6.66 0.00 6.66 0.00 4.86 5.94 4.86 5.94 3.74 6.26 3.74
                 6.26 4.86 12.93 4.86 12.93 3.96 13.25 3.96 13.25 4.86
                 15.40 4.86 15.40 4.80 15.80 4.80 15.80 4.86 19.20 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  17.84 3.89 15.75 3.89 15.75 4.16 13.64 4.16 13.64 3.53
                 13.57 3.53 13.57 3.18 12.42 3.18 12.42 2.86 13.57 2.86
                 13.57 1.22 13.89 1.22 13.89 3.21 13.96 3.21 13.96 3.84
                 15.43 3.84 15.43 3.57 17.52 3.57 17.52 2.34 17.84 2.34 ;
        POLYGON  13.25 2.47 12.93 2.47 12.93 2.28 11.03 2.28 11.03 4.54
                 10.71 4.54 10.71 2.28 10.27 1.84 10.27 1.22 10.59 1.22
                 10.59 1.70 10.85 1.96 13.25 1.96 ;
        RECT  11.49 3.96 12.49 4.28 ;
        RECT  11.09 1.22 12.39 1.54 ;
        POLYGON  10.39 3.90 9.33 3.90 9.33 3.58 10.07 3.58 10.07 2.60 9.65 2.18
                 7.51 2.18 7.29 2.40 7.29 2.58 6.97 2.58 6.97 2.26 7.37 1.86
                 9.79 1.86 10.39 2.46 ;
        RECT  7.37 4.22 10.33 4.54 ;
        RECT  7.13 1.22 9.77 1.54 ;
        POLYGON  9.51 2.82 8.55 2.82 7.95 3.42 7.09 3.42 7.09 3.90 6.77 3.90
                 6.77 3.42 6.33 3.42 6.33 2.32 3.88 2.32 3.88 2.00 6.33 2.00
                 6.33 1.66 6.45 1.66 6.45 1.22 6.77 1.22 6.77 1.99 6.65 1.99
                 6.65 3.10 7.81 3.10 8.41 2.50 9.51 2.50 ;
        RECT  4.41 3.46 5.45 3.78 ;
        RECT  4.00 1.22 5.37 1.54 ;
        POLYGON  5.09 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 5.09 4.22 ;
        POLYGON  4.03 3.90 3.30 3.90 3.30 3.04 0.80 3.04 0.80 2.66 1.12 2.66
                 1.12 2.72 2.92 2.72 2.92 2.00 3.30 1.62 3.30 1.22 3.62 1.22
                 3.62 1.76 3.24 2.14 3.24 2.72 3.62 2.72 3.62 3.58 4.03 3.58 ;
        RECT  1.82 1.22 2.92 1.54 ;
        RECT  1.82 3.58 2.92 3.90 ;
    END
END dffp_4

MACRO dffp_2
    CLASS CORE ;
    FOREIGN dffp_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.64 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.03 3.46 8.84 3.46 8.80 3.50 8.80 3.90 8.48 3.90 8.48 3.36
                 8.70 3.14 9.03 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.42 2.08 2.06 2.40 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.81 1.98 14.56 1.98 14.56 3.06 14.81 3.06 14.81 3.38
                 14.24 3.38 14.24 1.64 14.81 1.64 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.48 4.54 15.90 4.54 15.90 4.22 16.16 4.22 16.16 1.77
                 15.90 1.77 15.90 1.45 16.48 1.45 ;
        END
    END qb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 0.90 15.52 0.90 15.52 1.24 15.20 1.24 15.20 0.90
                 13.19 0.90 13.19 1.14 12.87 1.14 12.87 0.90 6.07 0.90
                 6.07 1.14 5.75 1.14 5.75 0.90 1.32 0.90 1.32 1.34 1.00 1.34
                 1.00 0.90 0.00 0.90 0.00 -0.90 16.64 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 6.66 0.00 6.66 0.00 4.86 5.94 4.86 5.94 3.74 6.26 3.74
                 6.26 4.86 12.93 4.86 12.93 3.96 13.25 3.96 13.25 4.86
                 16.64 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  15.70 3.84 15.45 3.84 15.45 4.54 13.57 4.54 13.57 3.18
                 12.59 3.18 12.59 2.86 13.57 2.86 13.57 1.22 13.89 1.22
                 13.89 4.22 15.13 4.22 15.13 3.52 15.38 3.52 15.38 2.14
                 15.70 2.14 ;
        POLYGON  13.25 2.47 12.93 2.47 12.93 2.28 11.03 2.28 11.03 4.54
                 10.71 4.54 10.71 2.28 10.27 1.84 10.27 1.22 10.59 1.22
                 10.59 1.70 10.85 1.96 13.25 1.96 ;
        RECT  11.49 3.96 12.49 4.28 ;
        RECT  11.09 1.22 12.39 1.54 ;
        POLYGON  10.39 3.90 9.33 3.90 9.33 3.58 10.07 3.58 10.07 2.60 9.65 2.18
                 7.51 2.18 7.29 2.40 7.29 2.58 6.97 2.58 6.97 2.26 7.37 1.86
                 9.79 1.86 10.39 2.46 ;
        RECT  7.37 4.22 10.33 4.54 ;
        RECT  7.13 1.22 9.77 1.54 ;
        POLYGON  9.51 2.82 8.55 2.82 7.95 3.42 7.09 3.42 7.09 3.90 6.77 3.90
                 6.77 3.42 6.33 3.42 6.33 2.32 3.88 2.32 3.88 2.00 6.33 2.00
                 6.33 1.66 6.45 1.66 6.45 1.22 6.77 1.22 6.77 1.99 6.65 1.99
                 6.65 3.10 7.81 3.10 8.41 2.50 9.51 2.50 ;
        RECT  4.41 3.46 5.45 3.78 ;
        RECT  4.00 1.22 5.37 1.54 ;
        POLYGON  5.09 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 5.09 4.22 ;
        POLYGON  4.03 3.90 3.30 3.90 3.30 3.04 0.80 3.04 0.80 2.66 1.12 2.66
                 1.12 2.72 2.92 2.72 2.92 2.00 3.30 1.62 3.30 1.22 3.62 1.22
                 3.62 1.76 3.24 2.14 3.24 2.72 3.62 2.72 3.62 3.58 4.03 3.58 ;
        RECT  1.82 1.22 2.92 1.54 ;
        RECT  1.82 3.58 2.92 3.90 ;
    END
END dffp_2

MACRO dffp_1
    CLASS CORE ;
    FOREIGN dffp_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.64 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.03 3.46 8.84 3.46 8.80 3.50 8.80 3.90 8.48 3.90 8.48 3.36
                 8.70 3.14 9.03 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.42 2.08 2.06 2.40 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.42  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.81 3.68 14.24 3.68 14.24 1.22 14.57 1.22 14.57 1.56
                 14.56 1.56 14.56 3.36 14.81 3.36 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.48 4.54 15.97 4.54 15.97 4.22 16.16 4.22 16.16 1.55
                 15.65 1.55 15.65 1.23 16.48 1.23 ;
        END
    END qb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 0.90 15.27 0.90 15.27 1.24 14.95 1.24 14.95 0.90
                 13.19 0.90 13.19 1.14 12.87 1.14 12.87 0.90 6.07 0.90
                 6.07 1.14 5.75 1.14 5.75 0.90 1.32 0.90 1.32 1.34 1.00 1.34
                 1.00 0.90 0.00 0.90 0.00 -0.90 16.64 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 6.66 0.00 6.66 0.00 4.86 5.94 4.86 5.94 3.74 6.26 3.74
                 6.26 4.86 12.93 4.86 12.93 3.96 13.25 3.96 13.25 4.86
                 16.64 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  15.45 4.54 13.57 4.54 13.57 3.18 12.59 3.18 12.59 2.86
                 13.57 2.86 13.57 1.22 13.89 1.22 13.89 4.22 15.13 4.22
                 15.13 2.46 15.11 2.46 15.11 2.14 15.45 2.14 ;
        POLYGON  13.25 2.47 12.93 2.47 12.93 2.28 11.03 2.28 11.03 4.54
                 10.71 4.54 10.71 2.28 10.27 1.84 10.27 1.22 10.59 1.22
                 10.59 1.70 10.85 1.96 13.25 1.96 ;
        RECT  11.49 3.96 12.49 4.28 ;
        RECT  11.09 1.22 12.39 1.54 ;
        POLYGON  10.39 3.90 9.33 3.90 9.33 3.58 10.07 3.58 10.07 2.60 9.65 2.18
                 7.51 2.18 7.29 2.40 7.29 2.58 6.97 2.58 6.97 2.26 7.37 1.86
                 9.79 1.86 10.39 2.46 ;
        RECT  7.37 4.22 10.33 4.54 ;
        RECT  7.13 1.22 9.77 1.54 ;
        POLYGON  9.51 2.82 8.55 2.82 7.95 3.42 7.09 3.42 7.09 3.90 6.77 3.90
                 6.77 3.42 6.33 3.42 6.33 2.32 3.88 2.32 3.88 2.00 6.33 2.00
                 6.33 1.66 6.45 1.66 6.45 1.22 6.77 1.22 6.77 1.99 6.65 1.99
                 6.65 3.10 7.81 3.10 8.41 2.50 9.51 2.50 ;
        RECT  4.41 3.46 5.45 3.78 ;
        RECT  4.00 1.22 5.37 1.54 ;
        POLYGON  5.09 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 5.09 4.22 ;
        POLYGON  4.03 3.90 3.30 3.90 3.30 3.04 0.80 3.04 0.80 2.66 1.12 2.66
                 1.12 2.72 2.92 2.72 2.92 2.00 3.30 1.62 3.30 1.22 3.62 1.22
                 3.62 1.76 3.24 2.14 3.24 2.72 3.62 2.72 3.62 3.58 4.03 3.58 ;
        RECT  1.82 1.22 2.92 1.54 ;
        RECT  1.82 3.58 2.92 3.90 ;
    END
END dffp_1

MACRO dffnsqb_4
    CLASS CORE ;
    FOREIGN dffnsqb_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.20 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.51  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.25 2.92 9.44 2.92 9.44 3.04 9.12 3.04 9.12 2.60 10.25 2.60 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.44 2.94 3.04 2.94 3.04 3.04 2.72 3.04 2.72 2.62 3.44 2.62 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  19.04 4.53 17.17 4.53 17.17 4.21 18.72 4.21 18.72 1.90
                 17.17 1.90 17.17 1.58 19.04 1.58 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.99  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.76 3.46 1.14 3.46 1.14 3.14 1.44 3.14 1.44 2.72 1.76 2.72 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  19.20 0.90 18.20 0.90 18.20 1.24 17.86 1.24 17.86 0.90
                 14.73 0.90 14.73 1.54 14.41 1.54 14.41 0.90 7.12 0.90
                 7.12 1.48 6.80 1.48 6.80 0.90 2.86 0.90 2.86 1.28 2.54 1.28
                 2.54 0.90 0.00 0.90 0.00 -0.90 19.20 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  19.20 6.66 0.00 6.66 0.00 4.86 2.54 4.86 2.54 4.60 2.86 4.60
                 2.86 4.86 7.36 4.86 7.36 3.74 7.68 3.74 7.68 4.86 9.75 4.86
                 9.75 4.36 10.07 4.36 10.07 4.86 13.37 4.86 13.37 4.60
                 13.69 4.60 13.69 4.86 15.51 4.86 15.51 3.96 15.83 3.96
                 15.83 4.86 19.20 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  18.19 3.89 16.39 3.89 16.39 3.18 15.49 3.18 15.49 3.64
                 14.07 3.64 14.07 3.32 15.17 3.32 15.17 2.86 16.39 2.86
                 16.39 1.88 16.49 1.88 16.49 1.22 16.81 1.22 16.81 2.20
                 16.71 2.20 16.71 3.57 17.87 3.57 17.87 2.34 18.19 2.34 ;
        RECT  15.11 1.22 16.11 1.54 ;
        POLYGON  16.07 2.47 15.75 2.47 15.75 2.28 12.23 2.28 12.23 4.54
                 11.91 4.54 11.91 2.02 11.77 1.88 11.77 1.22 12.09 1.22
                 12.09 1.74 12.31 1.96 16.07 1.96 ;
        RECT  12.69 3.96 15.07 4.28 ;
        RECT  12.47 1.22 14.03 1.54 ;
        POLYGON  11.53 4.04 9.89 4.04 9.89 3.68 9.37 3.68 9.37 4.32 9.05 4.32
                 9.05 3.36 10.21 3.36 10.21 3.72 11.53 3.72 ;
        POLYGON  11.51 3.40 10.53 3.40 10.53 3.08 11.19 3.08 11.19 2.34
                 11.03 2.18 8.08 2.18 8.08 1.86 11.17 1.86 11.51 2.20 ;
        RECT  8.72 1.22 11.39 1.54 ;
        POLYGON  8.51 4.48 8.19 4.48 8.19 2.82 5.88 2.82 5.88 3.06 5.56 3.06
                 5.56 2.50 7.44 2.50 7.44 1.22 8.38 1.22 8.38 1.54 7.76 1.54
                 7.76 2.50 8.51 2.50 ;
        RECT  5.83 3.46 6.87 3.78 ;
        POLYGON  6.51 4.54 3.18 4.54 3.18 4.28 2.16 4.28 2.16 4.54 0.46 4.54
                 0.46 1.22 0.78 1.22 0.78 4.22 1.84 4.22 1.84 3.96 3.50 3.96
                 3.50 4.22 6.51 4.22 ;
        RECT  5.42 1.22 6.42 1.54 ;
        POLYGON  5.45 3.90 4.72 3.90 4.72 2.18 2.49 2.18 2.49 2.38 2.17 2.38
                 2.17 1.86 4.72 1.86 4.72 1.22 5.04 1.22 5.04 3.58 5.45 3.58 ;
        RECT  3.24 1.22 4.34 1.54 ;
        RECT  3.24 3.32 4.34 3.64 ;
        RECT  1.16 1.22 2.16 1.54 ;
    END
END dffnsqb_4

MACRO dffnsqb_2
    CLASS CORE ;
    FOREIGN dffnsqb_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.56 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.51  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.25 2.92 9.44 2.92 9.44 3.04 9.12 3.04 9.12 2.60 10.25 2.60 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.44 2.94 3.04 2.94 3.04 3.04 2.72 3.04 2.72 2.62 3.44 2.62 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  18.40 4.32 17.87 4.32 17.87 4.00 18.08 4.00 18.08 1.55
                 17.87 1.55 17.87 1.23 18.40 1.23 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.99  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.76 3.46 1.14 3.46 1.14 3.14 1.44 3.14 1.44 2.72 1.76 2.72 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  18.56 0.90 17.49 0.90 17.49 1.54 17.17 1.54 17.17 0.90
                 14.73 0.90 14.73 1.54 14.41 1.54 14.41 0.90 7.12 0.90
                 7.12 1.48 6.80 1.48 6.80 0.90 2.86 0.90 2.86 1.28 2.54 1.28
                 2.54 0.90 0.00 0.90 0.00 -0.90 18.56 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  18.56 6.66 0.00 6.66 0.00 4.86 2.54 4.86 2.54 4.60 2.86 4.60
                 2.86 4.86 7.36 4.86 7.36 3.74 7.68 3.74 7.68 4.86 9.75 4.86
                 9.75 4.36 10.07 4.36 10.07 4.86 13.37 4.86 13.37 4.60
                 13.69 4.60 13.69 4.86 15.51 4.86 15.51 3.96 15.83 3.96
                 15.83 4.86 18.56 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  17.70 3.68 17.43 3.68 17.43 4.54 16.39 4.54 16.39 3.18
                 15.49 3.18 15.49 3.64 14.07 3.64 14.07 3.32 15.17 3.32
                 15.17 2.86 16.49 2.86 16.49 1.22 16.81 1.22 16.81 3.18
                 16.71 3.18 16.71 4.22 17.11 4.22 17.11 3.36 17.38 3.36
                 17.38 2.46 17.33 2.46 17.33 2.14 17.70 2.14 ;
        POLYGON  16.17 2.47 15.85 2.47 15.85 2.28 12.23 2.28 12.23 4.54
                 11.91 4.54 11.91 2.02 11.77 1.88 11.77 1.22 12.09 1.22
                 12.09 1.74 12.31 1.96 16.17 1.96 ;
        RECT  15.11 1.22 16.11 1.54 ;
        RECT  12.69 3.96 15.07 4.28 ;
        RECT  12.47 1.22 14.03 1.54 ;
        POLYGON  11.53 4.04 9.89 4.04 9.89 3.68 9.05 3.68 9.05 3.36 10.21 3.36
                 10.21 3.72 11.53 3.72 ;
        POLYGON  11.51 3.40 10.53 3.40 10.53 3.08 11.19 3.08 11.19 2.34
                 11.03 2.18 8.08 2.18 8.08 1.86 11.17 1.86 11.51 2.20 ;
        RECT  8.72 1.22 11.39 1.54 ;
        POLYGON  8.51 4.48 8.19 4.48 8.19 2.82 5.88 2.82 5.88 3.06 5.56 3.06
                 5.56 2.50 7.44 2.50 7.44 1.22 8.38 1.22 8.38 1.54 7.76 1.54
                 7.76 2.50 8.51 2.50 ;
        RECT  5.83 3.46 6.87 3.78 ;
        POLYGON  6.51 4.54 3.18 4.54 3.18 4.28 2.16 4.28 2.16 4.54 0.46 4.54
                 0.46 1.22 0.78 1.22 0.78 4.22 1.84 4.22 1.84 3.96 3.50 3.96
                 3.50 4.22 6.51 4.22 ;
        RECT  5.42 1.22 6.42 1.54 ;
        POLYGON  5.45 3.90 4.72 3.90 4.72 2.18 2.49 2.18 2.49 2.38 2.17 2.38
                 2.17 1.86 4.72 1.86 4.72 1.22 5.04 1.22 5.04 3.58 5.45 3.58 ;
        RECT  3.24 1.22 4.34 1.54 ;
        RECT  3.24 3.32 4.34 3.64 ;
        RECT  1.16 1.22 2.16 1.54 ;
    END
END dffnsqb_2

MACRO dffnsqb_1
    CLASS CORE ;
    FOREIGN dffnsqb_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.56 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.51  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.25 2.92 9.44 2.92 9.44 3.04 9.12 3.04 9.12 2.60 10.25 2.60 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.44 2.94 3.04 2.94 3.04 3.04 2.72 3.04 2.72 2.62 3.44 2.62 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  18.40 4.32 17.87 4.32 17.87 4.00 18.08 4.00 18.08 1.55
                 17.87 1.55 17.87 1.23 18.40 1.23 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.99  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.76 3.46 1.14 3.46 1.14 3.14 1.44 3.14 1.44 2.72 1.76 2.72 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  18.56 0.90 17.49 0.90 17.49 1.54 17.17 1.54 17.17 0.90
                 14.73 0.90 14.73 1.54 14.41 1.54 14.41 0.90 7.12 0.90
                 7.12 1.48 6.80 1.48 6.80 0.90 2.86 0.90 2.86 1.28 2.54 1.28
                 2.54 0.90 0.00 0.90 0.00 -0.90 18.56 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  18.56 6.66 0.00 6.66 0.00 4.86 2.54 4.86 2.54 4.60 2.86 4.60
                 2.86 4.86 7.36 4.86 7.36 3.74 7.68 3.74 7.68 4.86 9.75 4.86
                 9.75 4.36 10.07 4.36 10.07 4.86 13.37 4.86 13.37 4.60
                 13.69 4.60 13.69 4.86 15.51 4.86 15.51 3.96 15.83 3.96
                 15.83 4.86 18.56 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  17.70 3.68 17.43 3.68 17.43 4.54 16.39 4.54 16.39 3.18
                 15.49 3.18 15.49 3.64 14.07 3.64 14.07 3.32 15.17 3.32
                 15.17 2.86 16.49 2.86 16.49 1.22 16.81 1.22 16.81 3.18
                 16.71 3.18 16.71 4.22 17.11 4.22 17.11 3.36 17.38 3.36
                 17.38 2.46 17.33 2.46 17.33 2.14 17.70 2.14 ;
        POLYGON  16.17 2.47 15.85 2.47 15.85 2.28 12.23 2.28 12.23 4.54
                 11.91 4.54 11.91 2.02 11.77 1.88 11.77 1.22 12.09 1.22
                 12.09 1.74 12.31 1.96 16.17 1.96 ;
        RECT  15.11 1.22 16.11 1.54 ;
        RECT  12.69 3.96 15.07 4.28 ;
        RECT  12.47 1.22 14.03 1.54 ;
        POLYGON  11.53 4.04 9.89 4.04 9.89 3.68 9.05 3.68 9.05 3.36 10.21 3.36
                 10.21 3.72 11.53 3.72 ;
        POLYGON  11.51 3.40 10.53 3.40 10.53 3.08 11.19 3.08 11.19 2.34
                 11.03 2.18 8.08 2.18 8.08 1.86 11.17 1.86 11.51 2.20 ;
        RECT  8.72 1.22 11.39 1.54 ;
        POLYGON  8.51 4.48 8.19 4.48 8.19 2.82 5.88 2.82 5.88 3.06 5.56 3.06
                 5.56 2.50 7.44 2.50 7.44 1.22 8.38 1.22 8.38 1.54 7.76 1.54
                 7.76 2.50 8.51 2.50 ;
        RECT  5.83 3.46 6.87 3.78 ;
        POLYGON  6.51 4.54 3.18 4.54 3.18 4.28 2.16 4.28 2.16 4.54 0.46 4.54
                 0.46 1.22 0.78 1.22 0.78 4.22 1.84 4.22 1.84 3.96 3.50 3.96
                 3.50 4.22 6.51 4.22 ;
        RECT  5.42 1.22 6.42 1.54 ;
        POLYGON  5.45 3.90 4.72 3.90 4.72 2.18 2.49 2.18 2.49 2.38 2.17 2.38
                 2.17 1.86 4.72 1.86 4.72 1.22 5.04 1.22 5.04 3.58 5.45 3.58 ;
        RECT  3.24 1.22 4.34 1.54 ;
        RECT  3.24 3.32 4.34 3.64 ;
        RECT  1.16 1.22 2.16 1.54 ;
    END
END dffnsqb_1

MACRO dffnsq_4
    CLASS CORE ;
    FOREIGN dffnsq_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.20 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.51  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.25 2.92 9.44 2.92 9.44 3.04 9.12 3.04 9.12 2.60 10.25 2.60 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.44 2.94 3.04 2.94 3.04 3.04 2.72 3.04 2.72 2.62 3.44 2.62 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  19.04 3.04 18.89 3.04 18.89 4.54 18.57 4.54 18.57 3.04
                 17.49 3.04 17.49 4.54 17.17 4.54 17.17 1.22 17.49 1.22
                 17.49 2.72 18.57 2.72 18.57 1.22 18.89 1.22 18.89 2.72
                 19.04 2.72 ;
        END
    END q
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.99  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.76 3.46 1.14 3.46 1.14 3.14 1.44 3.14 1.44 2.72 1.76 2.72 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  19.20 0.90 18.19 0.90 18.19 1.54 17.87 1.54 17.87 0.90
                 14.73 0.90 14.73 1.54 14.41 1.54 14.41 0.90 7.12 0.90
                 7.12 1.48 6.80 1.48 6.80 0.90 2.86 0.90 2.86 1.28 2.54 1.28
                 2.54 0.90 0.00 0.90 0.00 -0.90 19.20 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  19.20 6.66 0.00 6.66 0.00 4.86 2.54 4.86 2.54 4.60 2.86 4.60
                 2.86 4.86 7.36 4.86 7.36 3.74 7.68 3.74 7.68 4.86 9.75 4.86
                 9.75 4.36 10.07 4.36 10.07 4.86 13.37 4.86 13.37 4.60
                 13.69 4.60 13.69 4.86 15.51 4.86 15.51 3.96 15.83 3.96
                 15.83 4.86 17.87 4.86 17.87 3.58 18.19 3.58 18.19 4.86
                 19.20 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  16.81 2.04 16.71 2.04 16.71 4.32 16.39 4.32 16.39 3.18
                 15.49 3.18 15.49 3.64 14.07 3.64 14.07 3.32 15.17 3.32
                 15.17 2.86 16.39 2.86 16.39 1.72 16.49 1.72 16.49 1.22
                 16.81 1.22 ;
        RECT  15.11 1.22 16.11 1.54 ;
        POLYGON  16.07 2.47 15.75 2.47 15.75 2.28 12.23 2.28 12.23 4.54
                 11.91 4.54 11.91 2.02 11.77 1.88 11.77 1.22 12.09 1.22
                 12.09 1.74 12.31 1.96 16.07 1.96 ;
        RECT  12.69 3.96 15.07 4.28 ;
        RECT  12.47 1.22 14.03 1.54 ;
        POLYGON  11.53 4.04 9.89 4.04 9.89 3.68 9.37 3.68 9.37 4.32 9.05 4.32
                 9.05 3.36 10.21 3.36 10.21 3.72 11.53 3.72 ;
        POLYGON  11.51 3.40 10.53 3.40 10.53 3.08 11.19 3.08 11.19 2.34
                 11.03 2.18 8.08 2.18 8.08 1.86 11.17 1.86 11.51 2.20 ;
        RECT  8.72 1.22 11.39 1.54 ;
        POLYGON  8.51 4.48 8.19 4.48 8.19 2.82 5.88 2.82 5.88 3.06 5.56 3.06
                 5.56 2.50 7.44 2.50 7.44 1.22 8.38 1.22 8.38 1.54 7.76 1.54
                 7.76 2.50 8.51 2.50 ;
        RECT  5.83 3.46 6.87 3.78 ;
        POLYGON  6.51 4.54 3.18 4.54 3.18 4.28 2.16 4.28 2.16 4.54 0.46 4.54
                 0.46 1.22 0.78 1.22 0.78 4.22 1.84 4.22 1.84 3.96 3.50 3.96
                 3.50 4.22 6.51 4.22 ;
        RECT  5.42 1.22 6.42 1.54 ;
        POLYGON  5.45 3.90 4.72 3.90 4.72 2.18 2.49 2.18 2.49 2.38 2.17 2.38
                 2.17 1.86 4.72 1.86 4.72 1.22 5.04 1.22 5.04 3.58 5.45 3.58 ;
        RECT  3.24 1.22 4.34 1.54 ;
        RECT  3.24 3.32 4.34 3.64 ;
        RECT  1.16 1.22 2.16 1.54 ;
    END
END dffnsq_4

MACRO dffnsq_2
    CLASS CORE ;
    FOREIGN dffnsq_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.56 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.51  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.25 2.92 9.44 2.92 9.44 3.04 9.12 3.04 9.12 2.60 10.25 2.60 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.44 2.94 3.04 2.94 3.04 3.04 2.72 3.04 2.72 2.62 3.44 2.62 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  18.40 3.04 18.19 3.04 18.19 4.32 17.87 4.32 17.87 1.64
                 18.19 1.64 18.19 2.72 18.40 2.72 ;
        END
    END q
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.99  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.76 3.46 1.14 3.46 1.14 3.14 1.44 3.14 1.44 2.72 1.76 2.72 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  18.56 0.90 17.49 0.90 17.49 1.97 17.17 1.97 17.17 0.90
                 14.73 0.90 14.73 1.54 14.41 1.54 14.41 0.90 7.12 0.90
                 7.12 1.48 6.80 1.48 6.80 0.90 2.86 0.90 2.86 1.28 2.54 1.28
                 2.54 0.90 0.00 0.90 0.00 -0.90 18.56 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  18.56 6.66 0.00 6.66 0.00 4.86 2.54 4.86 2.54 4.60 2.86 4.60
                 2.86 4.86 7.36 4.86 7.36 3.74 7.68 3.74 7.68 4.86 9.75 4.86
                 9.75 4.36 10.07 4.36 10.07 4.86 13.37 4.86 13.37 4.60
                 13.69 4.60 13.69 4.86 15.51 4.86 15.51 3.96 15.83 3.96
                 15.83 4.86 17.17 4.86 17.17 4.04 17.49 4.04 17.49 4.86
                 18.56 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  16.81 3.18 16.71 3.18 16.71 4.32 16.39 4.32 16.39 3.18
                 15.49 3.18 15.49 3.64 14.07 3.64 14.07 3.32 15.17 3.32
                 15.17 2.86 16.49 2.86 16.49 1.22 16.81 1.22 ;
        POLYGON  16.17 2.47 15.85 2.47 15.85 2.28 12.23 2.28 12.23 4.54
                 11.91 4.54 11.91 2.02 11.77 1.88 11.77 1.22 12.09 1.22
                 12.09 1.74 12.31 1.96 16.17 1.96 ;
        RECT  15.11 1.22 16.11 1.54 ;
        RECT  12.69 3.96 15.07 4.28 ;
        RECT  12.47 1.22 14.03 1.54 ;
        POLYGON  11.53 4.04 9.89 4.04 9.89 3.68 9.37 3.68 9.37 4.32 9.05 4.32
                 9.05 3.36 10.21 3.36 10.21 3.72 11.53 3.72 ;
        POLYGON  11.51 3.40 10.53 3.40 10.53 3.08 11.19 3.08 11.19 2.34
                 11.03 2.18 8.08 2.18 8.08 1.86 11.17 1.86 11.51 2.20 ;
        RECT  8.72 1.22 11.39 1.54 ;
        POLYGON  8.51 4.48 8.19 4.48 8.19 2.82 5.88 2.82 5.88 3.06 5.56 3.06
                 5.56 2.50 7.44 2.50 7.44 1.22 8.38 1.22 8.38 1.54 7.76 1.54
                 7.76 2.50 8.51 2.50 ;
        RECT  5.83 3.46 6.87 3.78 ;
        POLYGON  6.51 4.54 3.18 4.54 3.18 4.28 2.16 4.28 2.16 4.54 0.46 4.54
                 0.46 1.22 0.78 1.22 0.78 4.22 1.84 4.22 1.84 3.96 3.50 3.96
                 3.50 4.22 6.51 4.22 ;
        RECT  5.42 1.22 6.42 1.54 ;
        POLYGON  5.45 3.90 4.72 3.90 4.72 2.18 2.49 2.18 2.49 2.38 2.17 2.38
                 2.17 1.86 4.72 1.86 4.72 1.22 5.04 1.22 5.04 3.58 5.45 3.58 ;
        RECT  3.24 1.22 4.34 1.54 ;
        RECT  3.24 3.32 4.34 3.64 ;
        RECT  1.16 1.22 2.16 1.54 ;
    END
END dffnsq_2

MACRO dffnsq_1
    CLASS CORE ;
    FOREIGN dffnsq_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.56 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.51  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.25 2.92 9.44 2.92 9.44 3.04 9.12 3.04 9.12 2.60 10.25 2.60 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.44 2.94 3.04 2.94 3.04 3.04 2.72 3.04 2.72 2.62 3.44 2.62 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  18.40 3.04 18.19 3.04 18.19 4.08 17.87 4.08 17.87 1.22
                 18.19 1.22 18.19 2.72 18.40 2.72 ;
        END
    END q
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.99  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.76 3.46 1.14 3.46 1.14 3.14 1.44 3.14 1.44 2.72 1.76 2.72 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  18.56 0.90 17.49 0.90 17.49 1.55 17.17 1.55 17.17 0.90
                 14.73 0.90 14.73 1.54 14.41 1.54 14.41 0.90 7.12 0.90
                 7.12 1.48 6.80 1.48 6.80 0.90 2.86 0.90 2.86 1.28 2.54 1.28
                 2.54 0.90 0.00 0.90 0.00 -0.90 18.56 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  18.56 6.66 0.00 6.66 0.00 4.86 2.54 4.86 2.54 4.60 2.86 4.60
                 2.86 4.86 7.36 4.86 7.36 3.74 7.68 3.74 7.68 4.86 9.75 4.86
                 9.75 4.36 10.07 4.36 10.07 4.86 13.37 4.86 13.37 4.60
                 13.69 4.60 13.69 4.86 15.51 4.86 15.51 3.96 15.83 3.96
                 15.83 4.86 17.17 4.86 17.17 4.28 17.49 4.28 17.49 4.86
                 18.56 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  16.81 3.18 16.71 3.18 16.71 4.32 16.39 4.32 16.39 3.18
                 15.49 3.18 15.49 3.64 14.07 3.64 14.07 3.32 15.17 3.32
                 15.17 2.86 16.49 2.86 16.49 1.22 16.81 1.22 ;
        POLYGON  16.17 2.47 15.85 2.47 15.85 2.28 12.23 2.28 12.23 4.54
                 11.91 4.54 11.91 2.02 11.77 1.88 11.77 1.22 12.09 1.22
                 12.09 1.74 12.31 1.96 16.17 1.96 ;
        RECT  15.11 1.22 16.11 1.54 ;
        RECT  12.69 3.96 15.07 4.28 ;
        RECT  12.47 1.22 14.03 1.54 ;
        POLYGON  11.53 4.04 9.89 4.04 9.89 3.68 9.37 3.68 9.37 4.32 9.05 4.32
                 9.05 3.36 10.21 3.36 10.21 3.72 11.53 3.72 ;
        POLYGON  11.51 3.40 10.53 3.40 10.53 3.08 11.19 3.08 11.19 2.34
                 11.03 2.18 8.08 2.18 8.08 1.86 11.17 1.86 11.51 2.20 ;
        RECT  8.72 1.22 11.39 1.54 ;
        POLYGON  8.51 3.90 8.19 3.90 8.19 2.82 5.88 2.82 5.88 3.06 5.56 3.06
                 5.56 2.50 7.44 2.50 7.44 1.22 8.38 1.22 8.38 1.54 7.76 1.54
                 7.76 2.50 8.51 2.50 ;
        RECT  5.83 3.46 6.87 3.78 ;
        POLYGON  6.51 4.54 3.18 4.54 3.18 4.28 2.16 4.28 2.16 4.54 0.46 4.54
                 0.46 1.22 0.78 1.22 0.78 4.22 1.84 4.22 1.84 3.96 3.50 3.96
                 3.50 4.22 6.51 4.22 ;
        RECT  5.42 1.22 6.42 1.54 ;
        POLYGON  5.45 3.90 4.72 3.90 4.72 2.18 2.49 2.18 2.49 2.38 2.17 2.38
                 2.17 1.86 4.72 1.86 4.72 1.22 5.04 1.22 5.04 3.58 5.45 3.58 ;
        RECT  3.24 1.22 4.34 1.54 ;
        RECT  3.24 3.32 4.34 3.64 ;
        RECT  1.16 1.22 2.16 1.54 ;
    END
END dffnsq_1

MACRO dffns_4
    CLASS CORE ;
    FOREIGN dffns_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.76 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.51  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.25 2.92 9.44 2.92 9.44 3.04 9.12 3.04 9.12 2.60 10.25 2.60 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.44 2.94 3.04 2.94 3.04 3.04 2.72 3.04 2.72 2.62 3.44 2.62 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  19.27 3.25 17.07 3.25 17.07 2.93 18.72 2.93 18.72 2.71
                 18.95 2.71 18.95 1.54 17.39 1.54 17.39 1.22 19.27 1.22 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  21.60 4.53 19.63 4.53 19.63 4.21 21.28 4.21 21.28 1.90
                 19.63 1.90 19.63 1.58 21.60 1.58 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.99  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.76 3.46 1.14 3.46 1.14 3.14 1.44 3.14 1.44 2.72 1.76 2.72 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.76 0.90 20.66 0.90 20.66 1.24 20.32 1.24 20.32 0.90
                 14.73 0.90 14.73 1.54 14.41 1.54 14.41 0.90 7.12 0.90
                 7.12 1.48 6.80 1.48 6.80 0.90 2.86 0.90 2.86 1.28 2.54 1.28
                 2.54 0.90 0.00 0.90 0.00 -0.90 21.76 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.76 6.66 0.00 6.66 0.00 4.86 2.54 4.86 2.54 4.60 2.86 4.60
                 2.86 4.86 7.36 4.86 7.36 3.74 7.68 3.74 7.68 4.86 9.75 4.86
                 9.75 4.36 10.07 4.36 10.07 4.86 13.37 4.86 13.37 4.60
                 13.69 4.60 13.69 4.86 15.51 4.86 15.51 3.96 15.83 3.96
                 15.83 4.86 17.73 4.86 17.73 4.80 18.13 4.80 18.13 4.86
                 21.76 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.65 3.89 16.39 3.89 16.39 3.18 15.49 3.18 15.49 3.64
                 14.07 3.64 14.07 3.32 15.17 3.32 15.17 2.86 16.39 2.86
                 16.39 1.88 16.49 1.88 16.49 1.22 16.81 1.22 16.81 2.20
                 16.71 2.20 16.71 3.57 20.33 3.57 20.33 2.34 20.65 2.34 ;
        RECT  15.11 1.22 16.11 1.54 ;
        POLYGON  16.07 2.47 15.75 2.47 15.75 2.28 12.23 2.28 12.23 4.54
                 11.91 4.54 11.91 2.02 11.77 1.88 11.77 1.22 12.09 1.22
                 12.09 1.74 12.31 1.96 16.07 1.96 ;
        RECT  12.69 3.96 15.07 4.28 ;
        RECT  12.47 1.22 14.03 1.54 ;
        POLYGON  11.53 4.04 9.89 4.04 9.89 3.68 9.37 3.68 9.37 4.32 9.05 4.32
                 9.05 3.36 10.21 3.36 10.21 3.72 11.53 3.72 ;
        POLYGON  11.51 3.40 10.53 3.40 10.53 3.08 11.19 3.08 11.19 2.34
                 11.03 2.18 8.08 2.18 8.08 1.86 11.17 1.86 11.51 2.20 ;
        RECT  8.72 1.22 11.39 1.54 ;
        POLYGON  8.51 4.48 8.19 4.48 8.19 2.82 5.88 2.82 5.88 3.06 5.56 3.06
                 5.56 2.50 7.44 2.50 7.44 1.22 8.38 1.22 8.38 1.54 7.76 1.54
                 7.76 2.50 8.51 2.50 ;
        RECT  5.83 3.46 6.87 3.78 ;
        POLYGON  6.51 4.54 3.18 4.54 3.18 4.28 2.16 4.28 2.16 4.54 0.46 4.54
                 0.46 1.22 0.78 1.22 0.78 4.22 1.84 4.22 1.84 3.96 3.50 3.96
                 3.50 4.22 6.51 4.22 ;
        RECT  5.42 1.22 6.42 1.54 ;
        POLYGON  5.45 3.90 4.72 3.90 4.72 2.18 2.49 2.18 2.49 2.38 2.17 2.38
                 2.17 1.86 4.72 1.86 4.72 1.22 5.04 1.22 5.04 3.58 5.45 3.58 ;
        RECT  3.24 1.22 4.34 1.54 ;
        RECT  3.24 3.32 4.34 3.64 ;
        RECT  1.16 1.22 2.16 1.54 ;
    END
END dffns_4

MACRO dffns_2
    CLASS CORE ;
    FOREIGN dffns_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.20 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.51  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.25 2.92 9.44 2.92 9.44 3.04 9.12 3.04 9.12 2.60 10.25 2.60 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.44 2.94 3.04 2.94 3.04 3.04 2.72 3.04 2.72 2.62 3.44 2.62 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  17.76 3.04 17.49 3.04 17.49 3.75 17.17 3.75 17.17 1.22
                 17.49 1.22 17.49 2.72 17.76 2.72 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  19.04 4.32 18.57 4.32 18.57 4.00 18.72 4.00 18.72 1.55
                 18.57 1.55 18.57 1.23 19.04 1.23 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.99  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.76 3.46 1.14 3.46 1.14 3.14 1.44 3.14 1.44 2.72 1.76 2.72 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  19.20 0.90 18.19 0.90 18.19 1.40 17.87 1.40 17.87 0.90
                 14.73 0.90 14.73 1.54 14.41 1.54 14.41 0.90 7.12 0.90
                 7.12 1.48 6.80 1.48 6.80 0.90 2.86 0.90 2.86 1.28 2.54 1.28
                 2.54 0.90 0.00 0.90 0.00 -0.90 19.20 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  19.20 6.66 0.00 6.66 0.00 4.86 2.54 4.86 2.54 4.60 2.86 4.60
                 2.86 4.86 7.36 4.86 7.36 3.74 7.68 3.74 7.68 4.86 9.75 4.86
                 9.75 4.36 10.07 4.36 10.07 4.86 13.37 4.86 13.37 4.60
                 13.69 4.60 13.69 4.86 15.51 4.86 15.51 3.96 15.83 3.96
                 15.83 4.86 19.20 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  18.40 3.68 18.13 3.68 18.13 4.54 16.39 4.54 16.39 3.18
                 15.49 3.18 15.49 3.64 14.07 3.64 14.07 3.32 15.17 3.32
                 15.17 2.86 16.49 2.86 16.49 1.22 16.81 1.22 16.81 3.18
                 16.71 3.18 16.71 4.22 17.81 4.22 17.81 3.36 18.08 3.36
                 18.08 2.46 18.03 2.46 18.03 2.14 18.40 2.14 ;
        POLYGON  16.17 2.47 15.85 2.47 15.85 2.28 12.23 2.28 12.23 4.54
                 11.91 4.54 11.91 2.02 11.77 1.88 11.77 1.22 12.09 1.22
                 12.09 1.74 12.31 1.96 16.17 1.96 ;
        RECT  15.11 1.22 16.11 1.54 ;
        RECT  12.69 3.96 15.07 4.28 ;
        RECT  12.47 1.22 14.03 1.54 ;
        POLYGON  11.53 4.04 9.89 4.04 9.89 3.68 9.05 3.68 9.05 3.36 10.21 3.36
                 10.21 3.72 11.53 3.72 ;
        POLYGON  11.51 3.40 10.53 3.40 10.53 3.08 11.19 3.08 11.19 2.34
                 11.03 2.18 8.08 2.18 8.08 1.86 11.17 1.86 11.51 2.20 ;
        RECT  8.72 1.22 11.39 1.54 ;
        POLYGON  8.51 4.48 8.19 4.48 8.19 2.82 5.88 2.82 5.88 3.06 5.56 3.06
                 5.56 2.50 7.44 2.50 7.44 1.22 8.38 1.22 8.38 1.54 7.76 1.54
                 7.76 2.50 8.51 2.50 ;
        RECT  5.83 3.46 6.87 3.78 ;
        POLYGON  6.51 4.54 3.18 4.54 3.18 4.28 2.16 4.28 2.16 4.54 0.46 4.54
                 0.46 1.22 0.78 1.22 0.78 4.22 1.84 4.22 1.84 3.96 3.50 3.96
                 3.50 4.22 6.51 4.22 ;
        RECT  5.42 1.22 6.42 1.54 ;
        POLYGON  5.45 3.90 4.72 3.90 4.72 2.18 2.49 2.18 2.49 2.38 2.17 2.38
                 2.17 1.86 4.72 1.86 4.72 1.22 5.04 1.22 5.04 3.58 5.45 3.58 ;
        RECT  3.24 1.22 4.34 1.54 ;
        RECT  3.24 3.32 4.34 3.64 ;
        RECT  1.16 1.22 2.16 1.54 ;
    END
END dffns_2

MACRO dffns_1
    CLASS CORE ;
    FOREIGN dffns_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.20 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.51  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.25 2.92 9.44 2.92 9.44 3.04 9.12 3.04 9.12 2.60 10.25 2.60 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.44 2.94 3.04 2.94 3.04 3.04 2.72 3.04 2.72 2.62 3.44 2.62 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.21  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  17.76 3.04 17.49 3.04 17.49 3.90 17.17 3.90 17.17 1.22
                 17.49 1.22 17.49 2.72 17.76 2.72 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.21  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  19.04 4.32 18.57 4.32 18.57 4.00 18.72 4.00 18.72 1.55
                 18.57 1.55 18.57 1.23 19.04 1.23 ;
        END
    END qb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.99  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.76 3.46 1.14 3.46 1.14 3.14 1.44 3.14 1.44 2.72 1.76 2.72 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  19.20 0.90 18.19 0.90 18.19 1.54 17.87 1.54 17.87 0.90
                 14.73 0.90 14.73 1.54 14.41 1.54 14.41 0.90 7.12 0.90
                 7.12 1.48 6.80 1.48 6.80 0.90 2.86 0.90 2.86 1.28 2.54 1.28
                 2.54 0.90 0.00 0.90 0.00 -0.90 19.20 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  19.20 6.66 0.00 6.66 0.00 4.86 2.54 4.86 2.54 4.60 2.86 4.60
                 2.86 4.86 7.36 4.86 7.36 3.74 7.68 3.74 7.68 4.86 9.75 4.86
                 9.75 4.36 10.07 4.36 10.07 4.86 13.37 4.86 13.37 4.60
                 13.69 4.60 13.69 4.86 15.51 4.86 15.51 3.96 15.83 3.96
                 15.83 4.86 19.20 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  18.40 3.68 18.13 3.68 18.13 4.54 16.39 4.54 16.39 3.18
                 15.49 3.18 15.49 3.64 14.07 3.64 14.07 3.32 15.17 3.32
                 15.17 2.86 16.49 2.86 16.49 1.22 16.81 1.22 16.81 3.18
                 16.71 3.18 16.71 4.22 17.81 4.22 17.81 3.36 18.08 3.36
                 18.08 2.46 18.03 2.46 18.03 2.14 18.40 2.14 ;
        POLYGON  16.17 2.47 15.85 2.47 15.85 2.28 12.23 2.28 12.23 4.54
                 11.91 4.54 11.91 2.02 11.77 1.88 11.77 1.22 12.09 1.22
                 12.09 1.74 12.31 1.96 16.17 1.96 ;
        RECT  15.11 1.22 16.11 1.54 ;
        RECT  12.69 3.96 15.07 4.28 ;
        RECT  12.47 1.22 14.03 1.54 ;
        POLYGON  11.53 4.04 9.89 4.04 9.89 3.68 9.05 3.68 9.05 3.36 10.21 3.36
                 10.21 3.72 11.53 3.72 ;
        POLYGON  11.51 3.40 10.53 3.40 10.53 3.08 11.19 3.08 11.19 2.34
                 11.03 2.18 8.08 2.18 8.08 1.86 11.17 1.86 11.51 2.20 ;
        RECT  8.72 1.22 11.39 1.54 ;
        POLYGON  8.51 4.48 8.19 4.48 8.19 2.82 5.88 2.82 5.88 3.06 5.56 3.06
                 5.56 2.50 7.44 2.50 7.44 1.22 8.38 1.22 8.38 1.54 7.76 1.54
                 7.76 2.50 8.51 2.50 ;
        RECT  5.83 3.46 6.87 3.78 ;
        POLYGON  6.51 4.54 3.18 4.54 3.18 4.28 2.16 4.28 2.16 4.54 0.46 4.54
                 0.46 1.22 0.78 1.22 0.78 4.22 1.84 4.22 1.84 3.96 3.50 3.96
                 3.50 4.22 6.51 4.22 ;
        RECT  5.42 1.22 6.42 1.54 ;
        POLYGON  5.45 3.90 4.72 3.90 4.72 2.18 2.49 2.18 2.49 2.38 2.17 2.38
                 2.17 1.86 4.72 1.86 4.72 1.22 5.04 1.22 5.04 3.58 5.45 3.58 ;
        RECT  3.24 1.22 4.34 1.54 ;
        RECT  3.24 3.32 4.34 3.64 ;
        RECT  1.16 1.22 2.16 1.54 ;
    END
END dffns_1

MACRO dffnrsqb_4
    CLASS CORE ;
    FOREIGN dffnrsqb_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.64 2.72 11.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.72 4.64 3.04 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  22.24 3.04 21.88 3.04 21.88 4.54 21.56 4.54 21.56 3.53
                 20.48 3.53 20.48 4.54 20.16 4.54 20.16 3.21 21.56 3.21
                 21.56 1.59 20.16 1.59 20.16 1.27 21.88 1.27 21.88 2.72
                 22.24 2.72 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.12 0.52 3.04 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.28 2.50 3.68 3.06 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  22.40 0.90 19.80 0.90 19.80 1.54 19.48 1.54 19.48 0.90
                 16.64 0.90 16.64 1.58 16.32 1.58 16.32 0.90 4.20 0.90
                 4.20 1.54 3.88 1.54 3.88 0.90 0.00 0.90 0.00 -0.90 22.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  22.40 6.66 0.00 6.66 0.00 4.86 0.99 4.86 0.99 4.16 1.31 4.16
                 1.31 4.86 5.52 4.86 5.52 4.62 5.84 4.62 5.84 4.86 9.40 4.86
                 9.40 4.16 9.72 4.16 9.72 4.86 11.68 4.86 11.68 4.64 12.00 4.64
                 12.00 4.86 15.32 4.86 15.32 3.94 15.64 3.94 15.64 4.86
                 19.48 4.86 19.48 4.22 19.80 4.22 19.80 4.86 20.86 4.86
                 20.86 4.22 21.18 4.22 21.18 4.86 22.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  19.96 2.70 19.10 2.70 19.10 3.06 18.42 3.06 18.42 3.90
                 18.10 3.90 18.10 3.06 17.02 3.06 17.02 4.54 16.70 4.54
                 16.70 2.90 15.92 2.90 15.92 2.58 17.02 2.58 17.02 2.74
                 18.78 2.74 18.78 1.22 19.10 1.22 19.10 2.36 19.96 2.36 ;
        POLYGON  19.10 4.54 17.40 4.54 17.40 3.58 17.72 3.58 17.72 4.22
                 19.10 4.22 ;
        POLYGON  18.12 2.42 17.79 2.42 17.79 2.22 14.56 2.22 14.56 2.70
                 14.16 3.10 14.16 4.12 13.84 4.12 13.84 2.96 14.24 2.56
                 14.24 1.26 14.56 1.26 14.56 1.90 18.12 1.90 ;
        RECT  17.02 1.26 18.02 1.58 ;
        POLYGON  16.34 3.62 14.86 3.62 14.86 3.80 14.54 3.80 14.54 3.30
                 16.34 3.30 ;
        RECT  14.94 1.26 15.94 1.58 ;
        POLYGON  13.86 1.58 13.54 1.58 13.54 1.54 11.30 1.54 11.30 1.22
                 13.86 1.22 ;
        RECT  10.90 4.00 13.46 4.32 ;
        POLYGON  13.42 3.08 13.12 3.08 13.12 3.68 12.46 3.68 12.46 3.36
                 12.80 3.36 12.80 2.18 10.66 2.18 10.66 1.54 9.10 1.54
                 9.10 2.58 7.84 2.58 7.84 2.84 7.52 2.84 7.52 2.26 8.78 2.26
                 8.78 1.22 10.98 1.22 10.98 1.86 13.18 1.86 13.18 2.18
                 13.12 2.18 13.12 2.76 13.42 2.76 ;
        POLYGON  12.48 2.92 12.14 2.92 12.14 3.68 9.74 3.68 9.74 3.22 8.42 3.22
                 8.42 2.90 9.74 2.90 9.74 1.86 10.10 1.86 10.10 2.18 10.06 2.18
                 10.06 3.36 11.82 3.36 11.82 2.58 12.48 2.58 ;
        RECT  7.70 3.58 8.90 3.90 ;
        RECT  7.00 1.22 8.46 1.54 ;
        POLYGON  8.46 4.54 6.52 4.54 6.52 4.30 4.14 4.30 4.14 3.70 1.68 3.70
                 1.68 2.42 1.58 2.42 1.58 1.22 1.90 1.22 1.90 2.10 2.00 2.10
                 2.00 3.38 4.46 3.38 4.46 3.98 6.84 3.98 6.84 4.22 8.46 4.22 ;
        POLYGON  7.32 3.70 7.00 3.70 7.00 3.26 6.76 3.02 5.96 3.02 5.96 2.18
                 2.96 2.18 2.96 2.98 2.64 2.98 2.64 1.86 5.96 1.86 5.96 1.22
                 6.30 1.22 6.30 1.54 6.28 1.54 6.28 2.70 6.90 2.70 7.32 3.12 ;
        RECT  4.82 3.34 6.62 3.66 ;
        RECT  4.60 1.22 5.60 1.54 ;
        RECT  1.82 4.02 3.63 4.34 ;
        RECT  2.28 1.22 3.28 1.54 ;
        POLYGON  1.36 2.98 1.16 2.98 1.16 3.72 0.50 3.72 0.50 4.54 0.18 4.54
                 0.18 3.40 0.84 3.40 0.84 1.54 0.18 1.54 0.18 1.22 1.16 1.22
                 1.16 2.66 1.36 2.66 ;
    END
END dffnrsqb_4

MACRO dffnrsqb_2
    CLASS CORE ;
    FOREIGN dffnrsqb_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.64 2.72 11.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.72 4.64 3.04 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.96 4.06 20.42 4.06 20.42 3.74 20.64 3.74 20.64 1.54
                 20.42 1.54 20.42 1.22 20.96 1.22 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.12 0.52 3.04 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.28 2.50 3.68 3.06 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 0.90 19.86 0.90 19.86 1.54 19.54 1.54 19.54 0.90
                 16.64 0.90 16.64 1.58 16.32 1.58 16.32 0.90 4.20 0.90
                 4.20 1.54 3.88 1.54 3.88 0.90 0.00 0.90 0.00 -0.90 21.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 6.66 0.00 6.66 0.00 4.86 0.99 4.86 0.99 4.16 1.31 4.16
                 1.31 4.86 5.52 4.86 5.52 4.62 5.84 4.62 5.84 4.86 9.40 4.86
                 9.40 4.16 9.72 4.16 9.72 4.86 11.68 4.86 11.68 4.64 12.00 4.64
                 12.00 4.86 15.32 4.86 15.32 3.94 15.64 3.94 15.64 4.86
                 19.60 4.86 19.60 4.22 19.92 4.22 19.92 4.86 21.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.32 3.06 18.42 3.06 18.42 3.90 18.10 3.90 18.10 3.06
                 17.02 3.06 17.02 4.54 16.70 4.54 16.70 2.90 15.92 2.90
                 15.92 2.58 17.02 2.58 17.02 2.74 18.78 2.74 18.78 1.22
                 19.10 1.22 19.10 2.74 20.00 2.74 20.00 2.62 20.32 2.62 ;
        POLYGON  19.10 4.54 17.40 4.54 17.40 3.58 17.72 3.58 17.72 4.22
                 19.10 4.22 ;
        POLYGON  18.12 2.42 17.79 2.42 17.79 2.22 14.56 2.22 14.56 2.70
                 14.16 3.10 14.16 4.12 13.84 4.12 13.84 2.96 14.24 2.56
                 14.24 1.26 14.56 1.26 14.56 1.90 18.12 1.90 ;
        RECT  17.02 1.26 18.02 1.58 ;
        POLYGON  16.34 3.62 14.86 3.62 14.86 3.80 14.54 3.80 14.54 3.30
                 16.34 3.30 ;
        RECT  14.94 1.26 15.94 1.58 ;
        POLYGON  13.86 1.58 13.54 1.58 13.54 1.54 11.30 1.54 11.30 1.22
                 13.86 1.22 ;
        RECT  10.90 4.00 13.46 4.32 ;
        POLYGON  13.42 3.08 13.12 3.08 13.12 3.68 12.46 3.68 12.46 3.36
                 12.80 3.36 12.80 2.18 10.66 2.18 10.66 1.54 9.10 1.54
                 9.10 2.58 7.84 2.58 7.84 2.84 7.52 2.84 7.52 2.26 8.78 2.26
                 8.78 1.22 10.98 1.22 10.98 1.86 13.18 1.86 13.18 2.18
                 13.12 2.18 13.12 2.76 13.42 2.76 ;
        POLYGON  12.48 2.92 12.14 2.92 12.14 3.68 9.74 3.68 9.74 3.22 8.42 3.22
                 8.42 2.90 9.74 2.90 9.74 1.86 10.10 1.86 10.10 2.18 10.06 2.18
                 10.06 3.36 11.82 3.36 11.82 2.58 12.48 2.58 ;
        RECT  7.70 3.58 8.90 3.90 ;
        RECT  7.00 1.22 8.46 1.54 ;
        POLYGON  8.46 4.54 6.52 4.54 6.52 4.30 4.14 4.30 4.14 3.70 1.68 3.70
                 1.68 2.42 1.58 2.42 1.58 1.22 1.90 1.22 1.90 2.10 2.00 2.10
                 2.00 3.38 4.46 3.38 4.46 3.98 6.84 3.98 6.84 4.22 8.46 4.22 ;
        POLYGON  7.32 3.70 7.00 3.70 7.00 3.26 6.76 3.02 5.96 3.02 5.96 2.18
                 2.96 2.18 2.96 2.98 2.64 2.98 2.64 1.86 5.96 1.86 5.96 1.22
                 6.30 1.22 6.30 1.54 6.28 1.54 6.28 2.70 6.90 2.70 7.32 3.12 ;
        RECT  4.82 3.34 6.62 3.66 ;
        RECT  4.60 1.22 5.60 1.54 ;
        RECT  1.82 4.02 3.63 4.34 ;
        RECT  2.28 1.22 3.28 1.54 ;
        POLYGON  1.36 2.98 1.16 2.98 1.16 3.72 0.50 3.72 0.50 4.54 0.18 4.54
                 0.18 3.40 0.84 3.40 0.84 1.54 0.18 1.54 0.18 1.22 1.16 1.22
                 1.16 2.66 1.36 2.66 ;
    END
END dffnrsqb_2

MACRO dffnrsqb_1
    CLASS CORE ;
    FOREIGN dffnrsqb_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.64 2.72 11.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.72 4.64 3.04 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.96 4.38 20.18 4.38 20.18 4.05 20.64 4.05 20.64 1.55
                 20.18 1.55 20.18 1.22 20.96 1.22 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.12 0.52 3.04 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.28 2.50 3.68 3.06 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 0.90 19.80 0.90 19.80 1.54 19.48 1.54 19.48 0.90
                 16.64 0.90 16.64 1.58 16.32 1.58 16.32 0.90 4.20 0.90
                 4.20 1.54 3.88 1.54 3.88 0.90 0.00 0.90 0.00 -0.90 21.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 6.66 0.00 6.66 0.00 4.86 0.99 4.86 0.99 4.16 1.31 4.16
                 1.31 4.86 5.52 4.86 5.52 4.62 5.84 4.62 5.84 4.86 9.40 4.86
                 9.40 4.16 9.72 4.16 9.72 4.86 11.68 4.86 11.68 4.64 12.00 4.64
                 12.00 4.86 15.32 4.86 15.32 3.94 15.64 3.94 15.64 4.86
                 21.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.08 3.06 18.42 3.06 18.42 3.90 18.10 3.90 18.10 3.06
                 17.02 3.06 17.02 4.54 16.70 4.54 16.70 2.90 15.92 2.90
                 15.92 2.58 17.02 2.58 17.02 2.74 18.60 2.74 18.60 1.22
                 18.92 1.22 18.92 2.74 19.76 2.74 19.76 2.62 20.08 2.62 ;
        POLYGON  19.10 4.54 17.40 4.54 17.40 3.58 17.72 3.58 17.72 4.22
                 19.10 4.22 ;
        POLYGON  18.12 2.42 17.79 2.42 17.79 2.22 14.56 2.22 14.56 2.70
                 14.16 3.10 14.16 4.12 13.84 4.12 13.84 2.96 14.24 2.56
                 14.24 1.26 14.56 1.26 14.56 1.90 18.12 1.90 ;
        RECT  17.02 1.26 18.02 1.58 ;
        POLYGON  16.34 3.62 14.86 3.62 14.86 3.80 14.54 3.80 14.54 3.30
                 16.34 3.30 ;
        RECT  14.94 1.26 15.94 1.58 ;
        POLYGON  13.86 1.58 13.54 1.58 13.54 1.54 11.30 1.54 11.30 1.22
                 13.86 1.22 ;
        RECT  10.90 4.00 13.46 4.32 ;
        POLYGON  13.42 3.08 13.12 3.08 13.12 3.68 12.46 3.68 12.46 3.36
                 12.80 3.36 12.80 2.18 10.66 2.18 10.66 1.54 9.10 1.54
                 9.10 2.58 7.84 2.58 7.84 2.84 7.52 2.84 7.52 2.26 8.78 2.26
                 8.78 1.22 10.98 1.22 10.98 1.86 13.18 1.86 13.18 2.18
                 13.12 2.18 13.12 2.76 13.42 2.76 ;
        POLYGON  12.48 2.92 12.14 2.92 12.14 3.68 9.74 3.68 9.74 3.22 8.42 3.22
                 8.42 2.90 9.74 2.90 9.74 1.86 10.10 1.86 10.10 2.18 10.06 2.18
                 10.06 3.36 11.82 3.36 11.82 2.58 12.48 2.58 ;
        RECT  7.70 3.58 8.90 3.90 ;
        RECT  7.00 1.22 8.46 1.54 ;
        POLYGON  8.46 4.54 6.52 4.54 6.52 4.30 4.14 4.30 4.14 3.70 1.68 3.70
                 1.68 2.42 1.58 2.42 1.58 1.22 1.90 1.22 1.90 2.10 2.00 2.10
                 2.00 3.38 4.46 3.38 4.46 3.98 6.84 3.98 6.84 4.22 8.46 4.22 ;
        POLYGON  7.32 3.70 7.00 3.70 7.00 3.26 6.76 3.02 5.96 3.02 5.96 2.18
                 2.96 2.18 2.96 2.98 2.64 2.98 2.64 1.86 5.96 1.86 5.96 1.22
                 6.30 1.22 6.30 1.54 6.28 1.54 6.28 2.70 6.90 2.70 7.32 3.12 ;
        RECT  4.82 3.34 6.62 3.66 ;
        RECT  4.60 1.22 5.60 1.54 ;
        RECT  1.82 4.02 3.63 4.34 ;
        RECT  2.28 1.22 3.28 1.54 ;
        POLYGON  1.36 2.98 1.16 2.98 1.16 3.72 0.50 3.72 0.50 4.54 0.18 4.54
                 0.18 3.40 0.84 3.40 0.84 1.54 0.18 1.54 0.18 1.22 1.16 1.22
                 1.16 2.66 1.36 2.66 ;
    END
END dffnrsqb_1

MACRO dffnrsq_4
    CLASS CORE ;
    FOREIGN dffnrsq_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.04 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.64 2.72 11.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.72 4.64 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  22.88 3.04 22.82 3.04 22.82 4.54 22.50 4.54 22.50 3.04
                 21.42 3.04 21.42 4.54 21.10 4.54 21.10 2.72 22.50 2.72
                 22.50 1.59 21.10 1.59 21.10 1.27 22.82 1.27 22.82 2.72
                 22.88 2.72 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.12 0.52 3.04 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.28 2.50 3.68 3.06 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  23.04 0.90 19.86 0.90 19.86 1.54 19.54 1.54 19.54 0.90
                 16.64 0.90 16.64 1.58 16.32 1.58 16.32 0.90 4.20 0.90
                 4.20 1.54 3.88 1.54 3.88 0.90 0.00 0.90 0.00 -0.90 23.04 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  23.04 6.66 0.00 6.66 0.00 4.86 0.99 4.86 0.99 4.16 1.31 4.16
                 1.31 4.86 5.52 4.86 5.52 4.62 5.84 4.62 5.84 4.86 9.40 4.86
                 9.40 4.16 9.72 4.16 9.72 4.86 11.68 4.86 11.68 4.64 12.00 4.64
                 12.00 4.86 15.32 4.86 15.32 3.94 15.64 3.94 15.64 4.86
                 19.60 4.86 19.60 4.22 19.92 4.22 19.92 4.86 21.80 4.86
                 21.80 3.58 22.12 3.58 22.12 4.86 23.04 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.90 2.45 20.74 2.45 20.74 4.54 20.42 4.54 20.42 1.22
                 20.74 1.22 20.74 2.13 20.90 2.13 ;
        POLYGON  20.10 3.06 18.42 3.06 18.42 3.90 18.10 3.90 18.10 3.06
                 17.02 3.06 17.02 4.54 16.70 4.54 16.70 2.90 15.92 2.90
                 15.92 2.58 17.02 2.58 17.02 2.74 18.78 2.74 18.78 1.22
                 19.10 1.22 19.10 2.74 19.78 2.74 19.78 2.62 20.10 2.62 ;
        POLYGON  19.10 4.54 17.40 4.54 17.40 3.58 17.72 3.58 17.72 4.22
                 19.10 4.22 ;
        POLYGON  18.12 2.42 17.79 2.42 17.79 2.22 14.56 2.22 14.56 2.70
                 14.16 3.10 14.16 4.12 13.84 4.12 13.84 2.96 14.24 2.56
                 14.24 1.26 14.56 1.26 14.56 1.90 18.12 1.90 ;
        RECT  17.02 1.26 18.02 1.58 ;
        POLYGON  16.34 3.62 14.86 3.62 14.86 3.80 14.54 3.80 14.54 3.30
                 16.34 3.30 ;
        RECT  14.94 1.26 15.94 1.58 ;
        POLYGON  13.86 1.58 13.54 1.58 13.54 1.54 11.30 1.54 11.30 1.22
                 13.86 1.22 ;
        RECT  10.90 4.00 13.46 4.32 ;
        POLYGON  13.42 3.08 13.12 3.08 13.12 3.68 12.46 3.68 12.46 3.36
                 12.80 3.36 12.80 2.18 10.66 2.18 10.66 1.54 9.10 1.54
                 9.10 2.58 7.84 2.58 7.84 2.84 7.52 2.84 7.52 2.26 8.78 2.26
                 8.78 1.22 10.98 1.22 10.98 1.86 13.18 1.86 13.18 2.18
                 13.12 2.18 13.12 2.76 13.42 2.76 ;
        POLYGON  12.48 2.92 12.14 2.92 12.14 3.68 9.74 3.68 9.74 3.22 8.42 3.22
                 8.42 2.90 9.74 2.90 9.74 1.86 10.10 1.86 10.10 2.18 10.06 2.18
                 10.06 3.36 11.82 3.36 11.82 2.58 12.48 2.58 ;
        RECT  7.70 3.58 8.90 3.90 ;
        RECT  7.00 1.22 8.46 1.54 ;
        POLYGON  8.46 4.54 6.52 4.54 6.52 4.30 4.14 4.30 4.14 3.70 1.68 3.70
                 1.68 2.42 1.58 2.42 1.58 1.22 1.90 1.22 1.90 2.10 2.00 2.10
                 2.00 3.38 4.46 3.38 4.46 3.98 6.84 3.98 6.84 4.22 8.46 4.22 ;
        POLYGON  7.32 3.70 7.00 3.70 7.00 3.26 6.76 3.02 5.96 3.02 5.96 2.18
                 2.96 2.18 2.96 2.98 2.64 2.98 2.64 1.86 5.96 1.86 5.96 1.22
                 6.30 1.22 6.30 1.54 6.28 1.54 6.28 2.70 6.90 2.70 7.32 3.12 ;
        RECT  4.82 3.34 6.62 3.66 ;
        RECT  4.60 1.22 5.60 1.54 ;
        RECT  1.82 4.02 3.63 4.34 ;
        RECT  2.28 1.22 3.28 1.54 ;
        POLYGON  1.36 2.98 1.16 2.98 1.16 3.72 0.50 3.72 0.50 4.54 0.18 4.54
                 0.18 3.40 0.84 3.40 0.84 1.54 0.18 1.54 0.18 1.22 1.16 1.22
                 1.16 2.66 1.36 2.66 ;
    END
END dffnrsq_4

MACRO dffnrsq_2
    CLASS CORE ;
    FOREIGN dffnrsq_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.64 2.72 11.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.72 4.64 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  22.24 3.04 22.12 3.04 22.12 4.54 21.80 4.54 21.80 1.64
                 22.12 1.64 22.12 2.72 22.24 2.72 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.12 0.52 3.04 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.28 2.50 3.68 3.06 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  22.40 0.90 21.42 0.90 21.42 1.96 21.10 1.96 21.10 0.90
                 19.86 0.90 19.86 1.54 19.54 1.54 19.54 0.90 16.64 0.90
                 16.64 1.58 16.32 1.58 16.32 0.90 4.20 0.90 4.20 1.54 3.88 1.54
                 3.88 0.90 0.00 0.90 0.00 -0.90 22.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  22.40 6.66 0.00 6.66 0.00 4.86 0.99 4.86 0.99 4.16 1.31 4.16
                 1.31 4.86 5.52 4.86 5.52 4.62 5.84 4.62 5.84 4.86 9.40 4.86
                 9.40 4.16 9.72 4.16 9.72 4.86 11.68 4.86 11.68 4.64 12.00 4.64
                 12.00 4.86 15.32 4.86 15.32 3.94 15.64 3.94 15.64 4.86
                 19.60 4.86 19.60 4.22 19.92 4.22 19.92 4.86 21.10 4.86
                 21.10 4.22 21.42 4.22 21.42 4.86 22.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.92 2.86 20.74 2.86 20.74 4.06 20.42 4.06 20.42 1.22
                 20.74 1.22 20.74 2.54 20.92 2.54 ;
        POLYGON  20.10 3.06 18.42 3.06 18.42 3.90 18.10 3.90 18.10 3.06
                 17.02 3.06 17.02 4.54 16.70 4.54 16.70 2.90 15.92 2.90
                 15.92 2.58 17.02 2.58 17.02 2.74 18.78 2.74 18.78 1.22
                 19.10 1.22 19.10 2.74 19.78 2.74 19.78 2.62 20.10 2.62 ;
        POLYGON  19.10 4.54 17.40 4.54 17.40 3.58 17.72 3.58 17.72 4.22
                 19.10 4.22 ;
        POLYGON  18.12 2.42 17.79 2.42 17.79 2.22 14.56 2.22 14.56 2.70
                 14.16 3.10 14.16 4.12 13.84 4.12 13.84 2.96 14.24 2.56
                 14.24 1.26 14.56 1.26 14.56 1.90 18.12 1.90 ;
        RECT  17.02 1.26 18.02 1.58 ;
        POLYGON  16.34 3.62 14.86 3.62 14.86 3.80 14.54 3.80 14.54 3.30
                 16.34 3.30 ;
        RECT  14.94 1.26 15.94 1.58 ;
        POLYGON  13.86 1.58 13.54 1.58 13.54 1.54 11.30 1.54 11.30 1.22
                 13.86 1.22 ;
        RECT  10.90 4.00 13.46 4.32 ;
        POLYGON  13.42 3.08 13.12 3.08 13.12 3.68 12.46 3.68 12.46 3.36
                 12.80 3.36 12.80 2.18 10.66 2.18 10.66 1.54 9.10 1.54
                 9.10 2.58 7.84 2.58 7.84 2.84 7.52 2.84 7.52 2.26 8.78 2.26
                 8.78 1.22 10.98 1.22 10.98 1.86 13.18 1.86 13.18 2.18
                 13.12 2.18 13.12 2.76 13.42 2.76 ;
        POLYGON  12.48 2.92 12.14 2.92 12.14 3.68 9.74 3.68 9.74 3.22 8.42 3.22
                 8.42 2.90 9.74 2.90 9.74 1.86 10.10 1.86 10.10 2.18 10.06 2.18
                 10.06 3.36 11.82 3.36 11.82 2.58 12.48 2.58 ;
        RECT  7.70 3.58 8.90 3.90 ;
        RECT  7.00 1.22 8.46 1.54 ;
        POLYGON  8.46 4.54 6.52 4.54 6.52 4.30 4.14 4.30 4.14 3.70 1.68 3.70
                 1.68 2.42 1.58 2.42 1.58 1.22 1.90 1.22 1.90 2.10 2.00 2.10
                 2.00 3.38 4.46 3.38 4.46 3.98 6.84 3.98 6.84 4.22 8.46 4.22 ;
        POLYGON  7.32 3.70 7.00 3.70 7.00 3.26 6.76 3.02 5.96 3.02 5.96 2.18
                 2.96 2.18 2.96 2.98 2.64 2.98 2.64 1.86 5.96 1.86 5.96 1.22
                 6.30 1.22 6.30 1.54 6.28 1.54 6.28 2.70 6.90 2.70 7.32 3.12 ;
        RECT  4.82 3.34 6.62 3.66 ;
        RECT  4.60 1.22 5.60 1.54 ;
        RECT  1.82 4.02 3.63 4.34 ;
        RECT  2.28 1.22 3.28 1.54 ;
        POLYGON  1.36 2.98 1.16 2.98 1.16 3.72 0.50 3.72 0.50 4.54 0.18 4.54
                 0.18 3.40 0.84 3.40 0.84 1.54 0.18 1.54 0.18 1.22 1.16 1.22
                 1.16 2.66 1.36 2.66 ;
    END
END dffnrsq_2

MACRO dffnrsq_1
    CLASS CORE ;
    FOREIGN dffnrsq_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.64 2.72 11.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.72 4.64 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  22.24 3.04 22.12 3.04 22.12 4.54 21.80 4.54 21.80 1.22
                 22.12 1.22 22.12 2.72 22.24 2.72 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.12 0.52 3.04 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.28 2.50 3.68 3.06 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  22.40 0.90 21.42 0.90 21.42 1.54 21.10 1.54 21.10 0.90
                 19.91 0.90 19.91 1.54 19.59 1.54 19.59 0.90 16.64 0.90
                 16.64 1.58 16.32 1.58 16.32 0.90 4.20 0.90 4.20 1.54 3.88 1.54
                 3.88 0.90 0.00 0.90 0.00 -0.90 22.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  22.40 6.66 0.00 6.66 0.00 4.86 0.99 4.86 0.99 4.16 1.31 4.16
                 1.31 4.86 5.52 4.86 5.52 4.62 5.84 4.62 5.84 4.86 9.40 4.86
                 9.40 4.16 9.72 4.16 9.72 4.86 11.68 4.86 11.68 4.64 12.00 4.64
                 12.00 4.86 15.32 4.86 15.32 3.94 15.64 3.94 15.64 4.86
                 19.60 4.86 19.60 4.28 19.92 4.28 19.92 4.86 21.10 4.86
                 21.10 3.98 21.42 3.98 21.42 4.86 22.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.92 2.94 20.74 2.94 20.74 4.54 20.42 4.54 20.42 1.22
                 20.74 1.22 20.74 2.62 20.92 2.62 ;
        POLYGON  20.10 3.06 18.42 3.06 18.42 3.90 18.10 3.90 18.10 3.06
                 17.02 3.06 17.02 4.54 16.70 4.54 16.70 2.90 15.92 2.90
                 15.92 2.58 17.02 2.58 17.02 2.74 18.78 2.74 18.78 1.22
                 19.10 1.22 19.10 2.74 19.78 2.74 19.78 2.62 20.10 2.62 ;
        POLYGON  19.10 4.54 17.40 4.54 17.40 3.58 17.72 3.58 17.72 4.22
                 19.10 4.22 ;
        POLYGON  18.12 2.42 17.79 2.42 17.79 2.22 14.56 2.22 14.56 2.70
                 14.16 3.10 14.16 4.12 13.84 4.12 13.84 2.96 14.24 2.56
                 14.24 1.26 14.56 1.26 14.56 1.90 18.12 1.90 ;
        RECT  17.02 1.26 18.02 1.58 ;
        POLYGON  16.34 3.62 14.86 3.62 14.86 3.80 14.54 3.80 14.54 3.30
                 16.34 3.30 ;
        RECT  14.94 1.26 15.94 1.58 ;
        POLYGON  13.86 1.58 13.54 1.58 13.54 1.54 11.30 1.54 11.30 1.22
                 13.86 1.22 ;
        RECT  10.90 4.00 13.46 4.32 ;
        POLYGON  13.42 3.08 13.12 3.08 13.12 3.68 12.46 3.68 12.46 3.36
                 12.80 3.36 12.80 2.18 10.66 2.18 10.66 1.54 9.10 1.54
                 9.10 2.58 7.84 2.58 7.84 2.84 7.52 2.84 7.52 2.26 8.78 2.26
                 8.78 1.22 10.98 1.22 10.98 1.86 13.18 1.86 13.18 2.18
                 13.12 2.18 13.12 2.76 13.42 2.76 ;
        POLYGON  12.48 2.92 12.14 2.92 12.14 3.68 9.74 3.68 9.74 3.22 8.42 3.22
                 8.42 2.90 9.74 2.90 9.74 1.86 10.10 1.86 10.10 2.18 10.06 2.18
                 10.06 3.36 11.82 3.36 11.82 2.58 12.48 2.58 ;
        RECT  7.70 3.58 8.90 3.90 ;
        RECT  7.00 1.22 8.46 1.54 ;
        POLYGON  8.46 4.54 6.52 4.54 6.52 4.30 4.14 4.30 4.14 3.70 1.68 3.70
                 1.68 2.42 1.58 2.42 1.58 1.22 1.90 1.22 1.90 2.10 2.00 2.10
                 2.00 3.38 4.46 3.38 4.46 3.98 6.84 3.98 6.84 4.22 8.46 4.22 ;
        POLYGON  7.32 3.70 7.00 3.70 7.00 3.26 6.76 3.02 5.96 3.02 5.96 2.18
                 2.96 2.18 2.96 2.98 2.64 2.98 2.64 1.86 5.96 1.86 5.96 1.22
                 6.30 1.22 6.30 1.54 6.28 1.54 6.28 2.70 6.90 2.70 7.32 3.12 ;
        RECT  4.82 3.34 6.62 3.66 ;
        RECT  4.60 1.22 5.60 1.54 ;
        RECT  1.82 4.02 3.63 4.34 ;
        RECT  2.28 1.22 3.28 1.54 ;
        POLYGON  1.36 2.98 1.16 2.98 1.16 3.72 0.50 3.72 0.50 4.54 0.18 4.54
                 0.18 3.40 0.84 3.40 0.84 1.54 0.18 1.54 0.18 1.22 1.16 1.22
                 1.16 2.66 1.36 2.66 ;
    END
END dffnrsq_1

MACRO dffnrs_4
    CLASS CORE ;
    FOREIGN dffnrs_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 25.60 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.64 2.72 11.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.72 4.64 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  25.44 4.53 23.67 4.53 23.67 4.21 25.12 4.21 25.12 1.90
                 23.67 1.90 23.67 1.58 25.44 1.58 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  23.52 3.25 21.58 3.25 21.58 2.93 23.20 2.93 23.20 2.52
                 22.90 2.52 22.90 1.54 21.10 1.54 21.10 1.22 23.22 1.22
                 23.22 2.20 23.52 2.20 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.12 0.52 3.04 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.28 2.50 3.68 3.06 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  25.60 0.90 24.70 0.90 24.70 1.24 24.36 1.24 24.36 0.90
                 19.86 0.90 19.86 1.54 19.54 1.54 19.54 0.90 16.64 0.90
                 16.64 1.58 16.32 1.58 16.32 0.90 4.20 0.90 4.20 1.54 3.88 1.54
                 3.88 0.90 0.00 0.90 0.00 -0.90 25.60 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  25.60 6.66 0.00 6.66 0.00 4.86 0.99 4.86 0.99 4.16 1.31 4.16
                 1.31 4.86 5.52 4.86 5.52 4.62 5.84 4.62 5.84 4.86 9.40 4.86
                 9.40 4.16 9.72 4.16 9.72 4.86 11.68 4.86 11.68 4.64 12.00 4.64
                 12.00 4.86 15.32 4.86 15.32 3.94 15.64 3.94 15.64 4.86
                 19.60 4.86 19.60 4.41 19.92 4.41 19.92 4.86 22.25 4.86
                 22.25 4.80 22.65 4.80 22.65 4.86 25.60 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  24.69 3.89 22.60 3.89 22.60 4.09 20.42 4.09 20.42 1.22
                 20.74 1.22 20.74 3.77 22.28 3.77 22.28 3.57 24.37 3.57
                 24.37 2.34 24.69 2.34 ;
        POLYGON  20.10 3.06 18.42 3.06 18.42 3.90 18.10 3.90 18.10 3.06
                 17.02 3.06 17.02 4.54 16.70 4.54 16.70 2.90 15.92 2.90
                 15.92 2.58 17.02 2.58 17.02 2.74 18.78 2.74 18.78 1.22
                 19.10 1.22 19.10 2.74 19.78 2.74 19.78 2.62 20.10 2.62 ;
        POLYGON  19.10 4.54 17.40 4.54 17.40 3.58 17.72 3.58 17.72 4.22
                 19.10 4.22 ;
        POLYGON  18.12 2.42 17.79 2.42 17.79 2.22 14.56 2.22 14.56 2.70
                 14.16 3.10 14.16 4.12 13.84 4.12 13.84 2.96 14.24 2.56
                 14.24 1.26 14.56 1.26 14.56 1.90 18.12 1.90 ;
        RECT  17.02 1.26 18.02 1.58 ;
        POLYGON  16.34 3.62 14.86 3.62 14.86 3.80 14.54 3.80 14.54 3.30
                 16.34 3.30 ;
        RECT  14.94 1.26 15.94 1.58 ;
        POLYGON  13.86 1.58 13.54 1.58 13.54 1.54 11.30 1.54 11.30 1.22
                 13.86 1.22 ;
        RECT  10.90 4.00 13.46 4.32 ;
        POLYGON  13.42 3.08 13.12 3.08 13.12 3.68 12.46 3.68 12.46 3.36
                 12.80 3.36 12.80 2.18 10.66 2.18 10.66 1.54 9.10 1.54
                 9.10 2.58 7.84 2.58 7.84 2.84 7.52 2.84 7.52 2.26 8.78 2.26
                 8.78 1.22 10.98 1.22 10.98 1.86 13.18 1.86 13.18 2.18
                 13.12 2.18 13.12 2.76 13.42 2.76 ;
        POLYGON  12.48 2.92 12.14 2.92 12.14 3.68 9.74 3.68 9.74 3.22 8.42 3.22
                 8.42 2.90 9.74 2.90 9.74 1.86 10.10 1.86 10.10 2.18 10.06 2.18
                 10.06 3.36 11.82 3.36 11.82 2.58 12.48 2.58 ;
        RECT  7.70 3.58 8.90 3.90 ;
        RECT  7.00 1.22 8.46 1.54 ;
        POLYGON  8.46 4.54 6.52 4.54 6.52 4.30 4.14 4.30 4.14 3.70 1.68 3.70
                 1.68 2.42 1.58 2.42 1.58 1.22 1.90 1.22 1.90 2.10 2.00 2.10
                 2.00 3.38 4.46 3.38 4.46 3.98 6.84 3.98 6.84 4.22 8.46 4.22 ;
        POLYGON  7.32 3.70 7.00 3.70 7.00 3.26 6.76 3.02 5.96 3.02 5.96 2.18
                 2.96 2.18 2.96 2.98 2.64 2.98 2.64 1.86 5.96 1.86 5.96 1.22
                 6.30 1.22 6.30 1.54 6.28 1.54 6.28 2.70 6.90 2.70 7.32 3.12 ;
        RECT  4.82 3.34 6.62 3.66 ;
        RECT  4.60 1.22 5.60 1.54 ;
        RECT  1.82 4.02 3.63 4.34 ;
        RECT  2.28 1.22 3.28 1.54 ;
        POLYGON  1.36 2.98 1.16 2.98 1.16 3.72 0.50 3.72 0.50 4.54 0.18 4.54
                 0.18 3.40 0.84 3.40 0.84 1.54 0.18 1.54 0.18 1.22 1.16 1.22
                 1.16 2.66 1.36 2.66 ;
    END
END dffnrs_4

MACRO dffnrs_2
    CLASS CORE ;
    FOREIGN dffnrs_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.04 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.64 2.72 11.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.72 4.64 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  21.60 3.45 21.42 3.45 21.42 3.90 21.10 3.90 21.10 3.13
                 21.28 3.13 21.28 2.27 21.10 2.27 21.10 1.22 21.42 1.22
                 21.42 1.95 21.60 1.95 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  22.88 4.54 22.54 4.54 22.54 4.22 22.56 4.22 22.56 1.54
                 22.54 1.54 22.54 1.22 22.88 1.22 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.12 0.52 3.04 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.28 2.50 3.68 3.06 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  23.04 0.90 22.12 0.90 22.12 1.54 21.80 1.54 21.80 0.90
                 19.86 0.90 19.86 1.54 19.54 1.54 19.54 0.90 16.64 0.90
                 16.64 1.58 16.32 1.58 16.32 0.90 4.20 0.90 4.20 1.54 3.88 1.54
                 3.88 0.90 0.00 0.90 0.00 -0.90 23.04 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  23.04 6.66 0.00 6.66 0.00 4.86 0.99 4.86 0.99 4.16 1.31 4.16
                 1.31 4.86 5.52 4.86 5.52 4.62 5.84 4.62 5.84 4.86 9.40 4.86
                 9.40 4.16 9.72 4.16 9.72 4.86 11.68 4.86 11.68 4.64 12.00 4.64
                 12.00 4.86 15.32 4.86 15.32 3.94 15.64 3.94 15.64 4.86
                 23.04 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  22.24 4.09 21.79 4.54 19.78 4.54 19.78 3.06 18.42 3.06
                 18.42 3.90 18.10 3.90 18.10 3.06 17.02 3.06 17.02 4.54
                 16.70 4.54 16.70 2.90 15.92 2.90 15.92 2.58 17.02 2.58
                 17.02 2.74 18.78 2.74 18.78 1.22 19.10 1.22 19.10 2.74
                 19.78 2.74 19.78 2.62 20.10 2.62 20.10 4.22 21.65 4.22
                 21.92 3.95 21.92 2.38 22.24 2.38 ;
        POLYGON  20.92 2.86 20.74 2.86 20.74 3.90 20.42 3.90 20.42 1.22
                 20.74 1.22 20.74 2.54 20.92 2.54 ;
        POLYGON  19.10 4.54 17.40 4.54 17.40 3.58 17.72 3.58 17.72 4.22
                 19.10 4.22 ;
        POLYGON  18.12 2.42 17.79 2.42 17.79 2.22 14.56 2.22 14.56 2.70
                 14.16 3.10 14.16 4.12 13.84 4.12 13.84 2.96 14.24 2.56
                 14.24 1.26 14.56 1.26 14.56 1.90 18.12 1.90 ;
        RECT  17.02 1.26 18.02 1.58 ;
        POLYGON  16.34 3.62 14.86 3.62 14.86 3.80 14.54 3.80 14.54 3.30
                 16.34 3.30 ;
        RECT  14.94 1.26 15.94 1.58 ;
        POLYGON  13.86 1.58 13.54 1.58 13.54 1.54 11.30 1.54 11.30 1.22
                 13.86 1.22 ;
        RECT  10.90 4.00 13.46 4.32 ;
        POLYGON  13.42 3.08 13.12 3.08 13.12 3.68 12.46 3.68 12.46 3.36
                 12.80 3.36 12.80 2.18 10.66 2.18 10.66 1.54 9.10 1.54
                 9.10 2.58 7.84 2.58 7.84 2.84 7.52 2.84 7.52 2.26 8.78 2.26
                 8.78 1.22 10.98 1.22 10.98 1.86 13.18 1.86 13.18 2.18
                 13.12 2.18 13.12 2.76 13.42 2.76 ;
        POLYGON  12.48 2.92 12.14 2.92 12.14 3.68 9.74 3.68 9.74 3.22 8.42 3.22
                 8.42 2.90 9.74 2.90 9.74 1.86 10.10 1.86 10.10 2.18 10.06 2.18
                 10.06 3.36 11.82 3.36 11.82 2.58 12.48 2.58 ;
        RECT  7.70 3.58 8.90 3.90 ;
        RECT  7.00 1.22 8.46 1.54 ;
        POLYGON  8.46 4.54 6.52 4.54 6.52 4.30 4.14 4.30 4.14 3.70 1.68 3.70
                 1.68 2.42 1.58 2.42 1.58 1.22 1.90 1.22 1.90 2.10 2.00 2.10
                 2.00 3.38 4.46 3.38 4.46 3.98 6.84 3.98 6.84 4.22 8.46 4.22 ;
        POLYGON  7.32 3.70 7.00 3.70 7.00 3.26 6.76 3.02 5.96 3.02 5.96 2.18
                 2.96 2.18 2.96 2.98 2.64 2.98 2.64 1.86 5.96 1.86 5.96 1.22
                 6.30 1.22 6.30 1.54 6.28 1.54 6.28 2.70 6.90 2.70 7.32 3.12 ;
        RECT  4.82 3.34 6.62 3.66 ;
        RECT  4.60 1.22 5.60 1.54 ;
        RECT  2.28 1.22 3.28 1.54 ;
        POLYGON  1.36 2.98 1.16 2.98 1.16 3.72 0.50 3.72 0.50 4.54 0.18 4.54
                 0.18 3.40 0.84 3.40 0.84 1.54 0.18 1.54 0.18 1.22 1.16 1.22
                 1.16 2.66 1.36 2.66 ;
        RECT  1.82 4.02 3.63 4.34 ;
    END
END dffnrs_2

MACRO dffnrs_1
    CLASS CORE ;
    FOREIGN dffnrs_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.04 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.64 2.72 11.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.72 4.64 3.04 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.21  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  21.60 3.45 21.42 3.45 21.42 3.90 21.10 3.90 21.10 3.13
                 21.28 3.13 21.28 2.27 21.10 2.27 21.10 1.22 21.42 1.22
                 21.42 1.95 21.60 1.95 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.21  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  22.88 4.54 22.54 4.54 22.54 4.22 22.56 4.22 22.56 1.54
                 22.54 1.54 22.54 1.22 22.88 1.22 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.12 0.52 3.04 ;
        END
    END rb
    PIN sb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.28 2.50 3.68 3.06 ;
        END
    END sb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  23.04 0.90 22.12 0.90 22.12 1.54 21.80 1.54 21.80 0.90
                 19.86 0.90 19.86 1.54 19.54 1.54 19.54 0.90 16.64 0.90
                 16.64 1.58 16.32 1.58 16.32 0.90 4.20 0.90 4.20 1.54 3.88 1.54
                 3.88 0.90 0.00 0.90 0.00 -0.90 23.04 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  23.04 6.66 0.00 6.66 0.00 4.86 0.99 4.86 0.99 4.16 1.31 4.16
                 1.31 4.86 5.52 4.86 5.52 4.62 5.84 4.62 5.84 4.86 9.40 4.86
                 9.40 4.16 9.72 4.16 9.72 4.86 11.68 4.86 11.68 4.64 12.00 4.64
                 12.00 4.86 15.32 4.86 15.32 3.94 15.64 3.94 15.64 4.86
                 23.04 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  22.24 4.09 21.79 4.54 19.78 4.54 19.78 3.06 18.42 3.06
                 18.42 3.90 18.10 3.90 18.10 3.06 17.02 3.06 17.02 4.54
                 16.70 4.54 16.70 2.90 15.92 2.90 15.92 2.58 17.02 2.58
                 17.02 2.74 18.78 2.74 18.78 1.22 19.10 1.22 19.10 2.74
                 19.78 2.74 19.78 2.62 20.10 2.62 20.10 4.22 21.65 4.22
                 21.92 3.95 21.92 2.38 22.24 2.38 ;
        POLYGON  20.92 2.86 20.74 2.86 20.74 3.90 20.42 3.90 20.42 1.22
                 20.74 1.22 20.74 2.54 20.92 2.54 ;
        POLYGON  19.10 4.54 17.40 4.54 17.40 3.58 17.72 3.58 17.72 4.22
                 19.10 4.22 ;
        POLYGON  18.12 2.42 17.79 2.42 17.79 2.22 14.56 2.22 14.56 2.70
                 14.16 3.10 14.16 4.12 13.84 4.12 13.84 2.96 14.24 2.56
                 14.24 1.26 14.56 1.26 14.56 1.90 18.12 1.90 ;
        RECT  17.02 1.26 18.02 1.58 ;
        POLYGON  16.34 3.62 14.86 3.62 14.86 3.80 14.54 3.80 14.54 3.30
                 16.34 3.30 ;
        RECT  14.94 1.26 15.94 1.58 ;
        POLYGON  13.86 1.58 13.54 1.58 13.54 1.54 11.30 1.54 11.30 1.22
                 13.86 1.22 ;
        RECT  10.90 4.00 13.46 4.32 ;
        POLYGON  13.42 3.08 13.12 3.08 13.12 3.68 12.46 3.68 12.46 3.36
                 12.80 3.36 12.80 2.18 10.66 2.18 10.66 1.54 9.10 1.54
                 9.10 2.58 7.84 2.58 7.84 2.84 7.52 2.84 7.52 2.26 8.78 2.26
                 8.78 1.22 10.98 1.22 10.98 1.86 13.18 1.86 13.18 2.18
                 13.12 2.18 13.12 2.76 13.42 2.76 ;
        POLYGON  12.48 2.92 12.14 2.92 12.14 3.68 9.74 3.68 9.74 3.22 8.42 3.22
                 8.42 2.90 9.74 2.90 9.74 1.86 10.10 1.86 10.10 2.18 10.06 2.18
                 10.06 3.36 11.82 3.36 11.82 2.58 12.48 2.58 ;
        RECT  7.70 3.58 8.90 3.90 ;
        RECT  7.00 1.22 8.46 1.54 ;
        POLYGON  8.46 4.54 6.52 4.54 6.52 4.30 4.14 4.30 4.14 3.70 1.68 3.70
                 1.68 2.42 1.58 2.42 1.58 1.22 1.90 1.22 1.90 2.10 2.00 2.10
                 2.00 3.38 4.46 3.38 4.46 3.98 6.84 3.98 6.84 4.22 8.46 4.22 ;
        POLYGON  7.32 3.70 7.00 3.70 7.00 3.26 6.76 3.02 5.96 3.02 5.96 2.18
                 2.96 2.18 2.96 2.98 2.64 2.98 2.64 1.86 5.96 1.86 5.96 1.22
                 6.30 1.22 6.30 1.54 6.28 1.54 6.28 2.70 6.90 2.70 7.32 3.12 ;
        RECT  4.82 3.34 6.62 3.66 ;
        RECT  4.60 1.22 5.60 1.54 ;
        RECT  2.28 1.22 3.28 1.54 ;
        POLYGON  1.36 2.98 1.16 2.98 1.16 3.72 0.50 3.72 0.50 4.54 0.18 4.54
                 0.18 3.40 0.84 3.40 0.84 1.54 0.18 1.54 0.18 1.22 1.16 1.22
                 1.16 2.66 1.36 2.66 ;
        RECT  1.82 4.02 3.63 4.34 ;
    END
END dffnrs_1

MACRO dffnrqb_4
    CLASS CORE ;
    FOREIGN dffnrqb_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  7.84 2.72 8.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.08 3.04 2.44 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.96 4.53 19.08 4.53 19.08 4.21 20.64 4.21 20.64 1.90
                 19.08 1.90 19.08 1.58 20.96 1.58 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.22  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 2.08 2.44 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 0.90 20.11 0.90 20.11 1.24 19.77 1.24 19.77 0.90
                 17.78 0.90 17.78 1.54 17.46 1.54 17.46 0.90 8.36 0.90
                 8.36 1.54 8.04 1.54 8.04 0.90 1.20 0.90 1.20 1.54 0.88 1.54
                 0.88 0.90 0.00 0.90 0.00 -0.90 21.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 6.66 0.00 6.66 0.00 4.86 16.08 4.86 16.08 4.18
                 16.40 4.18 16.40 4.86 17.58 4.86 17.58 4.51 17.90 4.51
                 17.90 4.86 21.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.10 3.89 18.20 3.89 18.20 3.20 16.14 3.20 16.14 2.88
                 18.26 2.88 18.26 2.00 18.16 2.00 18.16 1.58 18.48 1.58
                 18.48 1.76 18.60 1.76 18.60 3.57 19.78 3.57 19.78 2.34
                 20.10 2.34 ;
        POLYGON  17.94 2.56 15.82 2.56 15.82 3.52 17.08 3.52 17.08 4.49
                 16.76 4.49 16.76 3.84 14.42 3.84 14.22 4.04 14.22 4.54
                 13.90 4.54 13.90 3.90 14.28 3.52 15.50 3.52 15.50 2.56
                 14.80 2.56 14.00 1.76 14.00 1.22 14.32 1.22 14.32 1.62
                 14.94 2.24 17.94 2.24 ;
        RECT  16.08 1.22 17.08 1.54 ;
        RECT  14.70 1.22 15.70 1.54 ;
        RECT  14.60 4.18 15.70 4.50 ;
        POLYGON  13.74 3.24 13.08 3.90 11.98 3.90 11.98 4.54 8.18 4.54
                 8.18 4.05 8.03 3.90 6.86 3.90 6.86 3.26 5.26 3.26 5.26 2.94
                 7.18 2.94 7.18 3.58 8.17 3.58 8.50 3.91 8.50 4.22 11.66 4.22
                 11.66 3.58 12.94 3.58 13.42 3.10 13.42 2.50 13.10 2.18
                 10.38 2.18 10.38 1.86 13.24 1.86 13.74 2.36 ;
        RECT  12.62 1.22 13.62 1.54 ;
        RECT  12.52 4.22 13.52 4.54 ;
        POLYGON  13.10 2.96 11.34 2.96 11.34 3.90 8.82 3.90 8.82 2.18 5.58 2.18
                 5.58 2.62 5.26 2.62 5.26 1.86 9.14 1.86 9.14 3.58 11.02 3.58
                 11.02 2.64 13.10 2.64 ;
        POLYGON  12.24 1.54 10.06 1.54 10.06 2.54 10.60 2.54 10.60 2.86
                 9.74 2.86 9.74 1.22 12.24 1.22 ;
        POLYGON  7.86 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 7.86 4.22 ;
        RECT  6.66 1.22 7.66 1.54 ;
        RECT  5.54 3.58 6.54 3.90 ;
        RECT  5.28 1.22 6.28 1.54 ;
        POLYGON  5.08 3.90 4.62 3.90 4.62 2.40 3.68 2.40 3.68 3.08 2.14 3.08
                 2.14 3.90 1.82 3.90 1.82 3.08 0.80 3.08 0.80 2.72 1.12 2.72
                 1.12 2.76 3.36 2.76 3.36 2.08 4.58 2.08 4.58 1.22 4.90 1.22
                 4.90 2.08 4.94 2.08 4.94 3.58 5.08 3.58 ;
        POLYGON  4.30 3.90 2.50 3.90 2.50 3.58 3.98 3.58 3.98 3.36 4.30 3.36 ;
        RECT  3.20 1.22 4.20 1.54 ;
        RECT  1.58 1.22 2.82 1.54 ;
    END
END dffnrqb_4

MACRO dffnrqb_2
    CLASS CORE ;
    FOREIGN dffnrqb_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 20.48 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  7.84 2.72 8.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.08 3.04 2.44 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.32 4.54 19.78 4.54 19.78 4.22 20.00 4.22 20.00 1.54
                 19.78 1.54 19.78 1.22 20.32 1.22 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.22  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 2.08 2.44 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 0.90 19.40 0.90 19.40 1.54 19.08 1.54 19.08 0.90
                 17.78 0.90 17.78 1.54 17.46 1.54 17.46 0.90 8.36 0.90
                 8.36 1.54 8.04 1.54 8.04 0.90 1.20 0.90 1.20 1.54 0.88 1.54
                 0.88 0.90 0.00 0.90 0.00 -0.90 20.48 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 6.66 0.00 6.66 0.00 4.86 16.08 4.86 16.08 4.12
                 16.40 4.12 16.40 4.86 17.58 4.86 17.58 4.56 17.90 4.56
                 17.90 4.86 20.48 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  19.44 2.44 18.60 2.44 18.60 4.22 18.72 4.22 18.72 4.54
                 18.28 4.54 18.28 3.16 16.14 3.16 16.14 2.84 18.28 2.84
                 18.28 1.54 18.16 1.54 18.16 1.22 18.60 1.22 18.60 2.12
                 19.44 2.12 ;
        POLYGON  17.96 2.52 15.82 2.52 15.82 3.48 17.08 3.48 17.08 4.54
                 16.76 4.54 16.76 3.80 14.46 3.80 14.22 4.04 14.22 4.54
                 13.90 4.54 13.90 3.90 14.32 3.48 15.50 3.48 15.50 2.52
                 14.76 2.52 14.00 1.76 14.00 1.22 14.32 1.22 14.32 1.62
                 14.90 2.20 17.96 2.20 ;
        RECT  16.08 1.22 17.08 1.54 ;
        RECT  14.70 1.22 15.70 1.54 ;
        RECT  14.60 4.12 15.70 4.44 ;
        POLYGON  13.74 3.24 13.08 3.90 11.98 3.90 11.98 4.54 8.18 4.54
                 8.18 4.05 8.03 3.90 6.86 3.90 6.86 3.26 5.26 3.26 5.26 2.94
                 7.18 2.94 7.18 3.58 8.17 3.58 8.50 3.91 8.50 4.22 11.66 4.22
                 11.66 3.58 12.94 3.58 13.42 3.10 13.42 2.50 13.10 2.18
                 10.38 2.18 10.38 1.86 13.24 1.86 13.74 2.36 ;
        RECT  12.62 1.22 13.62 1.54 ;
        RECT  12.52 4.22 13.52 4.54 ;
        POLYGON  13.10 2.96 11.34 2.96 11.34 3.90 8.82 3.90 8.82 2.18 5.58 2.18
                 5.58 2.62 5.26 2.62 5.26 1.86 9.14 1.86 9.14 3.58 11.02 3.58
                 11.02 2.64 13.10 2.64 ;
        POLYGON  12.24 1.54 10.06 1.54 10.06 2.54 10.60 2.54 10.60 2.86
                 9.74 2.86 9.74 1.22 12.24 1.22 ;
        POLYGON  7.86 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 7.86 4.22 ;
        RECT  6.66 1.22 7.66 1.54 ;
        RECT  5.54 3.58 6.54 3.90 ;
        RECT  5.28 1.22 6.28 1.54 ;
        POLYGON  5.08 3.90 4.62 3.90 4.62 2.40 3.68 2.40 3.68 3.08 2.14 3.08
                 2.14 3.90 1.82 3.90 1.82 3.08 0.80 3.08 0.80 2.72 1.12 2.72
                 1.12 2.76 3.36 2.76 3.36 2.08 4.58 2.08 4.58 1.22 4.90 1.22
                 4.90 2.08 4.94 2.08 4.94 3.58 5.08 3.58 ;
        POLYGON  4.30 3.90 2.50 3.90 2.50 3.58 3.98 3.58 3.98 3.36 4.30 3.36 ;
        RECT  3.20 1.22 4.20 1.54 ;
        RECT  1.58 1.22 2.82 1.54 ;
    END
END dffnrqb_2

MACRO dffnrqb_1
    CLASS CORE ;
    FOREIGN dffnrqb_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 20.48 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  7.84 2.72 8.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.08 3.04 2.44 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.32 4.54 19.78 4.54 19.78 4.22 20.00 4.22 20.00 1.54
                 19.78 1.54 19.78 1.22 20.32 1.22 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.22  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 2.08 2.44 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 0.90 19.40 0.90 19.40 1.54 19.08 1.54 19.08 0.90
                 17.78 0.90 17.78 1.54 17.46 1.54 17.46 0.90 8.36 0.90
                 8.36 1.54 8.04 1.54 8.04 0.90 1.20 0.90 1.20 1.54 0.88 1.54
                 0.88 0.90 0.00 0.90 0.00 -0.90 20.48 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 6.66 0.00 6.66 0.00 4.86 16.08 4.86 16.08 4.12
                 16.40 4.12 16.40 4.86 17.58 4.86 17.58 4.56 17.90 4.56
                 17.90 4.86 20.48 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  19.44 3.16 18.60 3.16 18.60 4.22 18.72 4.22 18.72 4.54
                 18.28 4.54 18.28 3.16 16.14 3.16 16.14 2.84 18.28 2.84
                 18.28 1.54 18.16 1.54 18.16 1.22 18.60 1.22 18.60 2.84
                 19.44 2.84 ;
        POLYGON  17.96 2.52 15.82 2.52 15.82 3.48 17.08 3.48 17.08 4.54
                 16.76 4.54 16.76 3.80 14.46 3.80 14.22 4.04 14.22 4.54
                 13.90 4.54 13.90 3.90 14.32 3.48 15.50 3.48 15.50 2.52
                 14.76 2.52 14.00 1.76 14.00 1.22 14.32 1.22 14.32 1.62
                 14.90 2.20 17.96 2.20 ;
        RECT  16.08 1.22 17.08 1.54 ;
        RECT  14.70 1.22 15.70 1.54 ;
        RECT  14.60 4.12 15.70 4.44 ;
        POLYGON  13.74 3.24 13.08 3.90 11.98 3.90 11.98 4.54 8.18 4.54
                 8.18 4.05 8.03 3.90 6.86 3.90 6.86 3.26 5.26 3.26 5.26 2.94
                 7.18 2.94 7.18 3.58 8.17 3.58 8.50 3.91 8.50 4.22 11.66 4.22
                 11.66 3.58 12.94 3.58 13.42 3.10 13.42 2.50 13.10 2.18
                 10.38 2.18 10.38 1.86 13.24 1.86 13.74 2.36 ;
        RECT  12.62 1.22 13.62 1.54 ;
        RECT  12.52 4.22 13.52 4.54 ;
        POLYGON  13.10 2.96 11.34 2.96 11.34 3.90 8.82 3.90 8.82 2.18 5.58 2.18
                 5.58 2.62 5.26 2.62 5.26 1.86 9.14 1.86 9.14 3.58 11.02 3.58
                 11.02 2.64 13.10 2.64 ;
        POLYGON  12.24 1.54 10.06 1.54 10.06 2.54 10.60 2.54 10.60 2.86
                 9.74 2.86 9.74 1.22 12.24 1.22 ;
        POLYGON  7.86 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 7.86 4.22 ;
        RECT  6.66 1.22 7.66 1.54 ;
        RECT  5.54 3.58 6.54 3.90 ;
        RECT  5.28 1.22 6.28 1.54 ;
        POLYGON  5.08 3.90 4.62 3.90 4.62 2.40 3.68 2.40 3.68 3.08 2.14 3.08
                 2.14 3.90 1.82 3.90 1.82 3.08 0.80 3.08 0.80 2.72 1.12 2.72
                 1.12 2.76 3.36 2.76 3.36 2.08 4.58 2.08 4.58 1.22 4.90 1.22
                 4.90 2.08 4.94 2.08 4.94 3.58 5.08 3.58 ;
        POLYGON  4.30 3.90 2.50 3.90 2.50 3.58 3.98 3.58 3.98 3.36 4.30 3.36 ;
        RECT  3.20 1.22 4.20 1.54 ;
        RECT  1.58 1.22 2.82 1.54 ;
    END
END dffnrqb_1

MACRO dffnrq_4
    CLASS CORE ;
    FOREIGN dffnrq_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  7.84 2.72 8.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.08 3.04 2.44 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.96 3.04 20.80 3.04 20.80 4.54 20.48 4.54 20.48 3.04
                 19.40 3.04 19.40 4.54 19.08 4.54 19.08 1.22 19.40 1.22
                 19.40 2.72 20.48 2.72 20.48 1.22 20.80 1.22 20.80 2.72
                 20.96 2.72 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.22  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 2.08 2.44 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 0.90 20.10 0.90 20.10 1.54 19.78 1.54 19.78 0.90
                 17.78 0.90 17.78 1.54 17.46 1.54 17.46 0.90 8.36 0.90
                 8.36 1.54 8.04 1.54 8.04 0.90 1.20 0.90 1.20 1.54 0.88 1.54
                 0.88 0.90 0.00 0.90 0.00 -0.90 21.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 6.66 0.00 6.66 0.00 4.86 16.08 4.86 16.08 4.12
                 16.40 4.12 16.40 4.86 17.58 4.86 17.58 4.56 17.90 4.56
                 17.90 4.86 19.78 4.86 19.78 3.58 20.10 3.58 20.10 4.86
                 21.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  18.72 4.54 18.28 4.54 18.28 3.16 16.14 3.16 16.14 2.84
                 18.28 2.84 18.28 1.54 18.16 1.54 18.16 1.22 18.60 1.22
                 18.60 4.22 18.72 4.22 ;
        POLYGON  17.96 2.52 15.82 2.52 15.82 3.48 17.08 3.48 17.08 4.54
                 16.76 4.54 16.76 3.80 14.46 3.80 14.22 4.04 14.22 4.54
                 13.90 4.54 13.90 3.90 14.32 3.48 15.50 3.48 15.50 2.52
                 14.76 2.52 14.00 1.76 14.00 1.22 14.32 1.22 14.32 1.62
                 14.90 2.20 17.96 2.20 ;
        RECT  16.08 1.22 17.08 1.54 ;
        RECT  14.70 1.22 15.70 1.54 ;
        RECT  14.60 4.12 15.70 4.44 ;
        RECT  12.62 1.22 13.62 1.54 ;
        RECT  12.52 4.22 13.52 4.54 ;
        POLYGON  13.10 2.96 11.34 2.96 11.34 3.90 8.82 3.90 8.82 2.18 5.58 2.18
                 5.58 2.62 5.26 2.62 5.26 1.86 9.14 1.86 9.14 3.58 11.02 3.58
                 11.02 2.64 13.10 2.64 ;
        POLYGON  12.24 1.54 10.06 1.54 10.06 2.54 10.60 2.54 10.60 2.86
                 9.74 2.86 9.74 1.22 12.24 1.22 ;
        POLYGON  7.86 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 7.86 4.22 ;
        RECT  6.66 1.22 7.66 1.54 ;
        RECT  5.54 3.58 6.54 3.90 ;
        RECT  5.28 1.22 6.28 1.54 ;
        POLYGON  5.08 3.90 4.62 3.90 4.62 2.40 3.68 2.40 3.68 3.08 2.14 3.08
                 2.14 3.90 1.82 3.90 1.82 3.08 0.80 3.08 0.80 2.72 1.12 2.72
                 1.12 2.76 3.36 2.76 3.36 2.08 4.58 2.08 4.58 1.22 4.90 1.22
                 4.90 2.08 4.94 2.08 4.94 3.58 5.08 3.58 ;
        POLYGON  4.30 3.90 2.50 3.90 2.50 3.58 3.98 3.58 3.98 3.36 4.30 3.36 ;
        RECT  3.20 1.22 4.20 1.54 ;
        RECT  1.58 1.22 2.82 1.54 ;
        POLYGON  13.74 3.24 13.08 3.90 11.98 3.90 11.98 4.54 8.18 4.54
                 8.18 4.05 8.03 3.90 6.86 3.90 6.86 3.26 5.26 3.26 5.26 2.94
                 7.18 2.94 7.18 3.58 8.17 3.58 8.50 3.91 8.50 4.22 11.66 4.22
                 11.66 3.58 12.94 3.58 13.42 3.10 13.42 2.50 13.10 2.18
                 10.38 2.18 10.38 1.86 13.24 1.86 13.74 2.36 ;
    END
END dffnrq_4

MACRO dffnrq_2
    CLASS CORE ;
    FOREIGN dffnrq_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 20.48 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  7.84 2.72 8.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.08 3.04 2.44 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.32 3.04 20.10 3.04 20.10 4.54 19.78 4.54 19.78 1.64
                 20.10 1.64 20.10 2.72 20.32 2.72 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.22  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 2.08 2.44 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 0.90 19.40 0.90 19.40 1.96 19.08 1.96 19.08 0.90
                 17.78 0.90 17.78 1.54 17.46 1.54 17.46 0.90 8.36 0.90
                 8.36 1.54 8.04 1.54 8.04 0.90 1.20 0.90 1.20 1.54 0.88 1.54
                 0.88 0.90 0.00 0.90 0.00 -0.90 20.48 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 6.66 0.00 6.66 0.00 4.86 16.08 4.86 16.08 4.12
                 16.40 4.12 16.40 4.86 17.54 4.86 17.54 3.62 17.86 3.62
                 17.86 4.86 19.08 4.86 19.08 4.22 19.40 4.22 19.40 4.86
                 20.48 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  18.72 4.54 18.28 4.54 18.28 3.16 16.14 3.16 16.14 2.84
                 18.28 2.84 18.28 1.54 18.16 1.54 18.16 1.22 18.60 1.22
                 18.60 4.22 18.72 4.22 ;
        POLYGON  17.96 2.52 15.82 2.52 15.82 3.48 17.08 3.48 17.08 4.54
                 16.76 4.54 16.76 3.80 14.46 3.80 14.22 4.04 14.22 4.54
                 13.90 4.54 13.90 3.90 14.32 3.48 15.50 3.48 15.50 2.52
                 14.76 2.52 14.00 1.76 14.00 1.22 14.32 1.22 14.32 1.62
                 14.90 2.20 17.96 2.20 ;
        RECT  16.08 1.22 17.08 1.54 ;
        RECT  14.70 1.22 15.70 1.54 ;
        RECT  14.60 4.12 15.70 4.44 ;
        POLYGON  13.74 3.24 13.08 3.90 11.98 3.90 11.98 4.54 8.18 4.54
                 8.18 4.05 8.03 3.90 6.86 3.90 6.86 3.26 5.26 3.26 5.26 2.94
                 7.18 2.94 7.18 3.58 8.17 3.58 8.50 3.91 8.50 4.22 11.66 4.22
                 11.66 3.58 12.94 3.58 13.42 3.10 13.42 2.50 13.10 2.18
                 10.38 2.18 10.38 1.86 13.24 1.86 13.74 2.36 ;
        RECT  12.62 1.22 13.62 1.54 ;
        RECT  12.52 4.22 13.52 4.54 ;
        POLYGON  13.10 2.96 11.34 2.96 11.34 3.90 8.82 3.90 8.82 2.18 5.58 2.18
                 5.58 2.62 5.26 2.62 5.26 1.86 9.14 1.86 9.14 3.58 11.02 3.58
                 11.02 2.64 13.10 2.64 ;
        POLYGON  12.24 1.54 10.06 1.54 10.06 2.54 10.60 2.54 10.60 2.86
                 9.74 2.86 9.74 1.22 12.24 1.22 ;
        POLYGON  7.86 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 7.86 4.22 ;
        RECT  6.66 1.22 7.66 1.54 ;
        RECT  5.54 3.58 6.54 3.90 ;
        RECT  5.28 1.22 6.28 1.54 ;
        POLYGON  5.08 3.90 4.62 3.90 4.62 2.40 3.68 2.40 3.68 3.08 2.14 3.08
                 2.14 3.90 1.82 3.90 1.82 3.08 0.80 3.08 0.80 2.72 1.12 2.72
                 1.12 2.76 3.36 2.76 3.36 2.08 4.58 2.08 4.58 1.22 4.90 1.22
                 4.90 2.08 4.94 2.08 4.94 3.58 5.08 3.58 ;
        POLYGON  4.30 3.90 2.50 3.90 2.50 3.58 3.98 3.58 3.98 3.36 4.30 3.36 ;
        RECT  3.20 1.22 4.20 1.54 ;
        RECT  1.58 1.22 2.82 1.54 ;
    END
END dffnrq_2

MACRO dffnrq_1
    CLASS CORE ;
    FOREIGN dffnrq_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 20.48 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  7.84 2.72 8.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.08 3.04 2.44 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.32 3.04 20.10 3.04 20.10 4.30 19.78 4.30 19.78 1.22
                 20.10 1.22 20.10 2.72 20.32 2.72 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.22  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 2.08 2.44 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 0.90 19.40 0.90 19.40 1.54 19.08 1.54 19.08 0.90
                 17.78 0.90 17.78 1.54 17.46 1.54 17.46 0.90 8.36 0.90
                 8.36 1.54 8.04 1.54 8.04 0.90 1.20 0.90 1.20 1.54 0.88 1.54
                 0.88 0.90 0.00 0.90 0.00 -0.90 20.48 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  20.48 6.66 0.00 6.66 0.00 4.86 16.08 4.86 16.08 4.12
                 16.40 4.12 16.40 4.86 17.58 4.86 17.58 4.56 17.90 4.56
                 17.90 4.86 19.08 4.86 19.08 4.06 19.40 4.06 19.40 4.86
                 20.48 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  18.72 4.54 18.28 4.54 18.28 3.16 16.14 3.16 16.14 2.84
                 18.28 2.84 18.28 1.54 18.16 1.54 18.16 1.22 18.60 1.22
                 18.60 4.22 18.72 4.22 ;
        POLYGON  17.96 2.52 15.82 2.52 15.82 3.48 17.08 3.48 17.08 4.54
                 16.76 4.54 16.76 3.80 14.46 3.80 14.22 4.04 14.22 4.54
                 13.90 4.54 13.90 3.90 14.32 3.48 15.50 3.48 15.50 2.52
                 14.76 2.52 14.00 1.76 14.00 1.22 14.32 1.22 14.32 1.62
                 14.90 2.20 17.96 2.20 ;
        RECT  16.08 1.22 17.08 1.54 ;
        RECT  14.70 1.22 15.70 1.54 ;
        RECT  14.60 4.12 15.70 4.44 ;
        POLYGON  13.74 3.24 13.08 3.90 11.98 3.90 11.98 4.54 8.18 4.54
                 8.18 4.05 8.03 3.90 6.86 3.90 6.86 3.26 5.26 3.26 5.26 2.94
                 7.18 2.94 7.18 3.58 8.17 3.58 8.50 3.91 8.50 4.22 11.66 4.22
                 11.66 3.58 12.94 3.58 13.42 3.10 13.42 2.50 13.10 2.18
                 10.38 2.18 10.38 1.86 13.24 1.86 13.74 2.36 ;
        RECT  12.62 1.22 13.62 1.54 ;
        RECT  12.52 4.22 13.52 4.54 ;
        POLYGON  13.10 2.96 11.34 2.96 11.34 3.90 8.82 3.90 8.82 2.18 5.58 2.18
                 5.58 2.62 5.26 2.62 5.26 1.86 9.14 1.86 9.14 3.58 11.02 3.58
                 11.02 2.64 13.10 2.64 ;
        POLYGON  12.24 1.54 10.06 1.54 10.06 2.54 10.60 2.54 10.60 2.86
                 9.74 2.86 9.74 1.22 12.24 1.22 ;
        POLYGON  7.86 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 7.86 4.22 ;
        RECT  6.66 1.22 7.66 1.54 ;
        RECT  5.54 3.58 6.54 3.90 ;
        RECT  5.28 1.22 6.28 1.54 ;
        POLYGON  5.08 3.90 4.62 3.90 4.62 2.40 3.68 2.40 3.68 3.08 2.14 3.08
                 2.14 3.90 1.82 3.90 1.82 3.08 0.80 3.08 0.80 2.72 1.12 2.72
                 1.12 2.76 3.36 2.76 3.36 2.08 4.58 2.08 4.58 1.22 4.90 1.22
                 4.90 2.08 4.94 2.08 4.94 3.58 5.08 3.58 ;
        POLYGON  4.30 3.90 2.50 3.90 2.50 3.58 3.98 3.58 3.98 3.36 4.30 3.36 ;
        RECT  3.20 1.22 4.20 1.54 ;
        RECT  1.58 1.22 2.82 1.54 ;
    END
END dffnrq_1

MACRO dffnr_4
    CLASS CORE ;
    FOREIGN dffnr_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  7.84 2.72 8.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.08 3.04 2.44 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  21.05 3.25 19.32 3.25 19.32 2.93 20.64 2.93 20.64 1.54
                 18.84 1.54 18.84 1.22 20.96 1.22 20.96 2.93 21.05 2.93 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  23.52 4.53 21.41 4.53 21.41 4.21 23.20 4.21 23.20 1.90
                 21.41 1.90 21.41 1.58 23.52 1.58 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.22  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 2.08 2.44 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  23.68 0.90 22.44 0.90 22.44 1.24 22.10 1.24 22.10 0.90
                 17.78 0.90 17.78 1.54 17.46 1.54 17.46 0.90 8.36 0.90
                 8.36 1.54 8.04 1.54 8.04 0.90 1.20 0.90 1.20 1.54 0.88 1.54
                 0.88 0.90 0.00 0.90 0.00 -0.90 23.68 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  23.68 6.66 0.00 6.66 0.00 4.86 16.08 4.86 16.08 4.18
                 16.40 4.18 16.40 4.86 17.58 4.86 17.58 4.56 17.90 4.56
                 17.90 4.86 19.99 4.86 19.99 4.80 20.39 4.80 20.39 4.86
                 23.68 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  22.43 3.89 20.34 3.89 20.34 4.00 18.20 4.00 18.20 3.20
                 16.14 3.20 16.14 2.88 18.26 2.88 18.26 2.00 18.16 2.00
                 18.16 1.58 18.48 1.58 18.48 1.76 18.60 1.76 18.60 3.68
                 20.02 3.68 20.02 3.57 22.11 3.57 22.11 2.34 22.43 2.34 ;
        POLYGON  17.94 2.56 15.82 2.56 15.82 3.52 17.08 3.52 17.08 4.54
                 16.76 4.54 16.76 3.84 14.42 3.84 14.22 4.04 14.22 4.54
                 13.90 4.54 13.90 3.90 14.28 3.52 15.50 3.52 15.50 2.56
                 14.80 2.56 14.00 1.76 14.00 1.22 14.32 1.22 14.32 1.62
                 14.94 2.24 17.94 2.24 ;
        RECT  16.08 1.22 17.08 1.54 ;
        RECT  14.70 1.22 15.70 1.54 ;
        RECT  14.60 4.18 15.70 4.50 ;
        POLYGON  13.74 3.24 13.08 3.90 11.98 3.90 11.98 4.54 8.18 4.54
                 8.18 4.05 8.03 3.90 6.86 3.90 6.86 3.26 5.26 3.26 5.26 2.94
                 7.18 2.94 7.18 3.58 8.17 3.58 8.50 3.91 8.50 4.22 11.66 4.22
                 11.66 3.58 12.94 3.58 13.42 3.10 13.42 2.50 13.10 2.18
                 10.38 2.18 10.38 1.86 13.24 1.86 13.74 2.36 ;
        RECT  12.62 1.22 13.62 1.54 ;
        RECT  12.52 4.22 13.52 4.54 ;
        POLYGON  13.10 2.96 11.34 2.96 11.34 3.90 8.82 3.90 8.82 2.18 5.58 2.18
                 5.58 2.62 5.26 2.62 5.26 1.86 9.14 1.86 9.14 3.58 11.02 3.58
                 11.02 2.64 13.10 2.64 ;
        POLYGON  12.24 1.54 10.06 1.54 10.06 2.54 10.60 2.54 10.60 2.86
                 9.74 2.86 9.74 1.22 12.24 1.22 ;
        POLYGON  7.86 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 7.86 4.22 ;
        RECT  6.66 1.22 7.66 1.54 ;
        RECT  5.54 3.58 6.54 3.90 ;
        RECT  5.28 1.22 6.28 1.54 ;
        POLYGON  5.08 3.90 4.62 3.90 4.62 2.40 3.68 2.40 3.68 3.08 2.14 3.08
                 2.14 3.90 1.82 3.90 1.82 3.08 0.80 3.08 0.80 2.72 1.12 2.72
                 1.12 2.76 3.36 2.76 3.36 2.08 4.58 2.08 4.58 1.22 4.90 1.22
                 4.90 2.08 4.94 2.08 4.94 3.58 5.08 3.58 ;
        POLYGON  4.30 3.90 2.50 3.90 2.50 3.58 3.98 3.58 3.98 3.36 4.30 3.36 ;
        RECT  3.20 1.22 4.20 1.54 ;
        RECT  1.58 1.22 2.82 1.54 ;
    END
END dffnr_4

MACRO dffnr_2
    CLASS CORE ;
    FOREIGN dffnr_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  7.84 2.72 8.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.08 3.04 2.44 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.99  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  19.68 2.40 19.36 2.40 19.36 3.08 19.40 3.08 19.40 3.40
                 19.04 3.40 19.04 1.22 19.40 1.22 19.40 1.54 19.36 1.54
                 19.36 2.08 19.68 2.08 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.96 4.54 20.62 4.54 20.62 4.22 20.64 4.22 20.64 1.54
                 20.62 1.54 20.62 1.22 20.96 1.22 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.22  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 2.08 2.44 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 0.90 20.18 0.90 20.18 1.19 19.86 1.19 19.86 0.90
                 17.78 0.90 17.78 1.54 17.46 1.54 17.46 0.90 8.36 0.90
                 8.36 1.54 8.04 1.54 8.04 0.90 1.20 0.90 1.20 1.54 0.88 1.54
                 0.88 0.90 0.00 0.90 0.00 -0.90 21.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 6.66 0.00 6.66 0.00 4.86 16.08 4.86 16.08 4.12
                 16.40 4.12 16.40 4.86 17.58 4.86 17.58 4.56 17.90 4.56
                 17.90 4.86 21.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.32 3.40 19.18 4.54 18.28 4.54 18.28 3.16 16.14 3.16
                 16.14 2.84 18.28 2.84 18.28 1.54 18.16 1.54 18.16 1.22
                 18.60 1.22 18.60 4.22 19.04 4.22 20.00 3.26 20.00 2.14
                 20.32 2.14 ;
        POLYGON  17.96 2.52 15.82 2.52 15.82 3.48 17.08 3.48 17.08 4.54
                 16.76 4.54 16.76 3.80 14.46 3.80 14.22 4.04 14.22 4.54
                 13.90 4.54 13.90 3.90 14.32 3.48 15.50 3.48 15.50 2.52
                 14.76 2.52 14.00 1.76 14.00 1.22 14.32 1.22 14.32 1.62
                 14.90 2.20 17.96 2.20 ;
        RECT  16.08 1.22 17.08 1.54 ;
        RECT  14.70 1.22 15.70 1.54 ;
        RECT  14.60 4.12 15.70 4.44 ;
        POLYGON  13.74 3.24 13.08 3.90 11.98 3.90 11.98 4.54 8.18 4.54
                 8.18 4.05 8.03 3.90 6.86 3.90 6.86 3.26 5.26 3.26 5.26 2.94
                 7.18 2.94 7.18 3.58 8.17 3.58 8.50 3.91 8.50 4.22 11.66 4.22
                 11.66 3.58 12.94 3.58 13.42 3.10 13.42 2.50 13.10 2.18
                 10.38 2.18 10.38 1.86 13.24 1.86 13.74 2.36 ;
        RECT  12.62 1.22 13.62 1.54 ;
        RECT  12.52 4.22 13.52 4.54 ;
        POLYGON  13.10 2.96 11.34 2.96 11.34 3.90 8.82 3.90 8.82 2.18 5.58 2.18
                 5.58 2.62 5.26 2.62 5.26 1.86 9.14 1.86 9.14 3.58 11.02 3.58
                 11.02 2.64 13.10 2.64 ;
        POLYGON  12.24 1.54 10.06 1.54 10.06 2.54 10.60 2.54 10.60 2.86
                 9.74 2.86 9.74 1.22 12.24 1.22 ;
        POLYGON  7.86 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 7.86 4.22 ;
        RECT  6.66 1.22 7.66 1.54 ;
        RECT  5.54 3.58 6.54 3.90 ;
        RECT  5.28 1.22 6.28 1.54 ;
        POLYGON  5.08 3.90 4.62 3.90 4.62 2.40 3.68 2.40 3.68 3.08 2.14 3.08
                 2.14 3.90 1.82 3.90 1.82 3.08 0.80 3.08 0.80 2.72 1.12 2.72
                 1.12 2.76 3.36 2.76 3.36 2.08 4.58 2.08 4.58 1.22 4.90 1.22
                 4.90 2.08 4.94 2.08 4.94 3.58 5.08 3.58 ;
        POLYGON  4.30 3.90 2.50 3.90 2.50 3.58 3.98 3.58 3.98 3.36 4.30 3.36 ;
        RECT  3.20 1.22 4.20 1.54 ;
        RECT  1.58 1.22 2.82 1.54 ;
    END
END dffnr_2

MACRO dffnr_1
    CLASS CORE ;
    FOREIGN dffnr_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  7.84 2.72 8.50 3.04 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.08 3.04 2.44 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.51  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  19.68 3.04 19.36 3.04 19.36 3.36 19.40 3.36 19.40 3.68
                 19.04 3.68 19.04 1.22 19.40 1.22 19.40 1.54 19.36 1.54
                 19.36 2.72 19.68 2.72 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.96 4.54 20.62 4.54 20.62 4.22 20.64 4.22 20.64 1.54
                 20.62 1.54 20.62 1.22 20.96 1.22 ;
        END
    END qb
    PIN rb
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.22  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.08 2.08 2.44 ;
        END
    END rb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 0.90 20.18 0.90 20.18 1.54 19.86 1.54 19.86 0.90
                 17.78 0.90 17.78 1.54 17.46 1.54 17.46 0.90 8.36 0.90
                 8.36 1.54 8.04 1.54 8.04 0.90 1.20 0.90 1.20 1.54 0.88 1.54
                 0.88 0.90 0.00 0.90 0.00 -0.90 21.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  21.12 6.66 0.00 6.66 0.00 4.86 16.08 4.86 16.08 4.12
                 16.40 4.12 16.40 4.86 17.58 4.86 17.58 4.56 17.90 4.56
                 17.90 4.86 21.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  20.32 3.68 19.46 4.54 18.28 4.54 18.28 3.16 16.14 3.16
                 16.14 2.84 18.28 2.84 18.28 1.54 18.16 1.54 18.16 1.22
                 18.60 1.22 18.60 4.22 19.32 4.22 20.00 3.54 20.00 2.46
                 19.96 2.46 19.96 2.14 20.32 2.14 ;
        POLYGON  17.96 2.52 15.82 2.52 15.82 3.48 17.08 3.48 17.08 4.54
                 16.76 4.54 16.76 3.80 14.46 3.80 14.22 4.04 14.22 4.54
                 13.90 4.54 13.90 3.90 14.32 3.48 15.50 3.48 15.50 2.52
                 14.76 2.52 14.00 1.76 14.00 1.22 14.32 1.22 14.32 1.62
                 14.90 2.20 17.96 2.20 ;
        RECT  16.08 1.22 17.08 1.54 ;
        RECT  14.70 1.22 15.70 1.54 ;
        RECT  14.60 4.12 15.70 4.44 ;
        POLYGON  13.74 3.24 13.08 3.90 11.98 3.90 11.98 4.54 8.18 4.54
                 8.18 4.05 8.03 3.90 6.86 3.90 6.86 3.26 5.26 3.26 5.26 2.94
                 7.18 2.94 7.18 3.58 8.17 3.58 8.50 3.91 8.50 4.22 11.66 4.22
                 11.66 3.58 12.94 3.58 13.42 3.10 13.42 2.50 13.10 2.18
                 10.38 2.18 10.38 1.86 13.24 1.86 13.74 2.36 ;
        RECT  12.62 1.22 13.62 1.54 ;
        RECT  12.52 4.22 13.52 4.54 ;
        POLYGON  13.10 2.96 11.34 2.96 11.34 3.90 8.82 3.90 8.82 2.18 5.58 2.18
                 5.58 2.62 5.26 2.62 5.26 1.86 9.14 1.86 9.14 3.58 11.02 3.58
                 11.02 2.64 13.10 2.64 ;
        POLYGON  12.24 1.54 10.06 1.54 10.06 2.54 10.60 2.54 10.60 2.86
                 9.74 2.86 9.74 1.22 12.24 1.22 ;
        POLYGON  7.86 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 7.86 4.22 ;
        RECT  6.66 1.22 7.66 1.54 ;
        RECT  5.54 3.58 6.54 3.90 ;
        RECT  5.28 1.22 6.28 1.54 ;
        POLYGON  5.08 3.90 4.62 3.90 4.62 2.40 3.68 2.40 3.68 3.08 2.14 3.08
                 2.14 3.90 1.82 3.90 1.82 3.08 0.80 3.08 0.80 2.72 1.12 2.72
                 1.12 2.76 3.36 2.76 3.36 2.08 4.58 2.08 4.58 1.22 4.90 1.22
                 4.90 2.08 4.94 2.08 4.94 3.58 5.08 3.58 ;
        POLYGON  4.30 3.90 2.50 3.90 2.50 3.58 3.98 3.58 3.98 3.36 4.30 3.36 ;
        RECT  3.20 1.22 4.20 1.54 ;
        RECT  1.58 1.22 2.82 1.54 ;
    END
END dffnr_1

MACRO dffnqb_4
    CLASS CORE ;
    FOREIGN dffnqb_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.64 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.03 3.46 8.16 3.46 8.16 3.68 7.84 3.68 7.84 3.14 9.03 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.42 2.08 2.30 2.40 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.48 4.54 14.49 4.54 14.49 4.22 16.16 4.22 16.16 1.91
                 14.49 1.91 14.49 1.59 16.48 1.59 ;
        END
    END qb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 0.90 15.51 0.90 15.51 1.24 15.19 1.24 15.19 0.90
                 13.03 0.90 13.03 1.14 12.71 1.14 12.71 0.90 5.70 0.90
                 5.70 1.48 5.38 1.48 5.38 0.90 1.32 0.90 1.32 1.34 1.00 1.34
                 1.00 0.90 0.00 0.90 0.00 -0.90 16.64 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 6.66 0.00 6.66 0.00 4.86 5.94 4.86 5.94 3.74 6.26 3.74
                 6.26 4.86 12.93 4.86 12.93 4.26 13.25 4.26 13.25 4.86
                 16.64 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  15.51 3.34 15.08 3.34 15.08 3.90 13.41 3.90 13.41 3.18
                 12.59 3.18 12.59 2.86 13.41 2.86 13.41 1.22 13.73 1.22
                 13.73 3.58 14.76 3.58 14.76 3.02 15.19 3.02 15.19 2.35
                 15.51 2.35 ;
        POLYGON  13.09 2.47 12.77 2.47 12.77 2.28 11.03 2.28 11.03 4.54
                 10.71 4.54 10.71 2.28 10.27 1.84 10.27 1.22 10.59 1.22
                 10.59 1.70 10.85 1.96 13.09 1.96 ;
        RECT  11.49 3.96 12.49 4.28 ;
        RECT  11.09 1.22 12.23 1.54 ;
        RECT  7.37 4.22 10.33 4.54 ;
        POLYGON  10.17 3.90 9.33 3.90 9.33 3.58 9.85 3.58 9.85 2.34 9.69 2.18
                 6.66 2.18 6.66 1.86 9.83 1.86 10.17 2.20 ;
        RECT  7.13 1.22 9.77 1.54 ;
        POLYGON  9.53 2.86 9.21 2.86 9.21 2.82 7.09 2.82 7.09 3.90 6.77 3.90
                 6.77 2.82 4.46 2.82 4.46 3.06 4.14 3.06 4.14 2.50 6.02 2.50
                 6.02 1.22 6.40 1.22 6.40 1.54 6.34 1.54 6.34 2.50 9.53 2.50 ;
        RECT  4.41 3.46 5.45 3.78 ;
        POLYGON  5.09 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 5.09 4.22 ;
        RECT  4.00 1.22 5.00 1.54 ;
        POLYGON  4.03 3.90 3.24 3.90 3.24 3.04 0.80 3.04 0.80 2.66 1.12 2.66
                 1.12 2.72 3.30 2.72 3.30 1.22 3.62 1.22 3.62 3.04 3.56 3.04
                 3.56 3.58 4.03 3.58 ;
        RECT  1.82 1.22 2.92 1.54 ;
        RECT  1.82 3.58 2.92 3.90 ;
    END
END dffnqb_4

MACRO dffnqb_2
    CLASS CORE ;
    FOREIGN dffnqb_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.00 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.03 3.46 8.16 3.46 8.16 3.68 7.84 3.68 7.84 3.14 9.03 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.42 2.08 2.30 2.40 ;
        END
    END d
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  15.84 4.44 15.19 4.44 15.19 4.12 15.52 4.12 15.52 1.96
                 15.19 1.96 15.19 1.64 15.84 1.64 ;
        END
    END qb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 0.90 14.81 0.90 14.81 1.24 14.49 1.24 14.49 0.90
                 13.19 0.90 13.19 1.14 12.87 1.14 12.87 0.90 5.70 0.90
                 5.70 1.48 5.38 1.48 5.38 0.90 1.32 0.90 1.32 1.34 1.00 1.34
                 1.00 0.90 0.00 0.90 0.00 -0.90 16.00 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 6.66 0.00 6.66 0.00 4.86 5.94 4.86 5.94 3.74 6.26 3.74
                 6.26 4.86 12.93 4.86 12.93 3.96 13.25 3.96 13.25 4.86
                 16.00 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  14.97 2.68 14.75 2.68 14.75 4.54 13.57 4.54 13.57 3.18
                 12.59 3.18 12.59 2.86 13.57 2.86 13.57 1.22 13.89 1.22
                 13.89 4.22 14.43 4.22 14.43 2.36 14.97 2.36 ;
        POLYGON  13.25 2.47 12.93 2.47 12.93 2.28 11.03 2.28 11.03 4.54
                 10.71 4.54 10.71 2.28 10.27 1.84 10.27 1.22 10.59 1.22
                 10.59 1.70 10.85 1.96 13.25 1.96 ;
        RECT  11.49 3.96 12.49 4.28 ;
        RECT  11.09 1.22 12.39 1.54 ;
        RECT  7.37 4.22 10.33 4.54 ;
        POLYGON  10.17 3.90 9.33 3.90 9.33 3.58 9.85 3.58 9.85 2.34 9.69 2.18
                 6.66 2.18 6.66 1.86 9.83 1.86 10.17 2.20 ;
        RECT  7.13 1.22 9.77 1.54 ;
        POLYGON  9.53 2.86 9.21 2.86 9.21 2.82 7.09 2.82 7.09 3.90 6.77 3.90
                 6.77 2.82 4.46 2.82 4.46 3.06 4.14 3.06 4.14 2.50 6.02 2.50
                 6.02 1.22 6.40 1.22 6.40 1.54 6.34 1.54 6.34 2.50 9.53 2.50 ;
        RECT  4.41 3.46 5.45 3.78 ;
        POLYGON  5.09 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 5.09 4.22 ;
        RECT  4.00 1.22 5.00 1.54 ;
        POLYGON  4.03 3.90 3.24 3.90 3.24 3.04 0.80 3.04 0.80 2.66 1.12 2.66
                 1.12 2.72 3.30 2.72 3.30 1.22 3.62 1.22 3.62 3.04 3.56 3.04
                 3.56 3.58 4.03 3.58 ;
        RECT  1.82 1.22 2.92 1.54 ;
        RECT  1.82 3.58 2.92 3.90 ;
    END
END dffnqb_2

MACRO dffnqb_1
    CLASS CORE ;
    FOREIGN dffnqb_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.00 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  15.84 4.08 15.19 4.08 15.19 3.76 15.52 3.76 15.52 1.54
                 14.95 1.54 14.95 1.22 15.84 1.22 ;
        END
    END qb
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.03 3.46 8.16 3.46 8.16 3.68 7.84 3.68 7.84 3.14 9.03 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.42 2.08 2.30 2.40 ;
        END
    END d
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 0.90 14.57 0.90 14.57 1.24 14.25 1.24 14.25 0.90
                 13.19 0.90 13.19 1.14 12.87 1.14 12.87 0.90 5.70 0.90
                 5.70 1.48 5.38 1.48 5.38 0.90 1.32 0.90 1.32 1.34 1.00 1.34
                 1.00 0.90 0.00 0.90 0.00 -0.90 16.00 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 6.66 0.00 6.66 0.00 4.86 5.94 4.86 5.94 3.74 6.26 3.74
                 6.26 4.86 12.93 4.86 12.93 3.96 13.25 3.96 13.25 4.86
                 16.00 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  14.73 4.54 13.57 4.54 13.57 3.18 12.59 3.18 12.59 2.86
                 13.57 2.86 13.57 1.22 13.89 1.22 13.89 4.22 14.41 4.22
                 14.41 2.14 14.73 2.14 ;
        POLYGON  13.25 2.47 12.93 2.47 12.93 2.28 11.03 2.28 11.03 4.54
                 10.71 4.54 10.71 2.28 10.27 1.84 10.27 1.22 10.59 1.22
                 10.59 1.70 10.85 1.96 13.25 1.96 ;
        RECT  11.49 3.96 12.49 4.28 ;
        RECT  11.09 1.22 12.39 1.54 ;
        RECT  7.37 4.22 10.33 4.54 ;
        POLYGON  10.17 3.90 9.33 3.90 9.33 3.58 9.85 3.58 9.85 2.34 9.69 2.18
                 6.66 2.18 6.66 1.86 9.83 1.86 10.17 2.20 ;
        RECT  7.13 1.22 9.77 1.54 ;
        POLYGON  9.53 2.86 9.21 2.86 9.21 2.82 7.09 2.82 7.09 3.90 6.77 3.90
                 6.77 2.82 4.46 2.82 4.46 3.06 4.14 3.06 4.14 2.50 6.02 2.50
                 6.02 1.22 6.40 1.22 6.40 1.54 6.34 1.54 6.34 2.50 9.53 2.50 ;
        RECT  4.41 3.46 5.45 3.78 ;
        POLYGON  5.09 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 5.09 4.22 ;
        RECT  4.00 1.22 5.00 1.54 ;
        POLYGON  4.03 3.90 3.24 3.90 3.24 3.04 0.80 3.04 0.80 2.66 1.12 2.66
                 1.12 2.72 3.30 2.72 3.30 1.22 3.62 1.22 3.62 3.04 3.56 3.04
                 3.56 3.58 4.03 3.58 ;
        RECT  1.82 1.22 2.92 1.54 ;
        RECT  1.82 3.58 2.92 3.90 ;
    END
END dffnqb_1

MACRO dffnq_4
    CLASS CORE ;
    FOREIGN dffnq_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.64 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.03 3.46 8.16 3.46 8.16 3.68 7.84 3.68 7.84 3.14 9.03 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.42 2.08 2.30 2.40 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.21 4.54 15.89 4.54 15.89 3.04 14.81 3.04 14.81 4.54
                 14.49 4.54 14.49 3.04 14.24 3.04 14.24 2.72 14.25 2.72
                 14.25 1.22 14.57 1.22 14.57 2.72 15.65 2.72 15.65 1.22
                 15.97 1.22 15.97 2.72 16.21 2.72 ;
        END
    END q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 0.90 15.27 0.90 15.27 1.54 14.95 1.54 14.95 0.90
                 13.19 0.90 13.19 1.14 12.87 1.14 12.87 0.90 5.70 0.90
                 5.70 1.48 5.38 1.48 5.38 0.90 1.32 0.90 1.32 1.34 1.00 1.34
                 1.00 0.90 0.00 0.90 0.00 -0.90 16.64 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 6.66 0.00 6.66 0.00 4.86 5.94 4.86 5.94 3.74 6.26 3.74
                 6.26 4.86 12.93 4.86 12.93 3.96 13.25 3.96 13.25 4.86
                 15.19 4.86 15.19 3.70 15.51 3.70 15.51 4.86 16.64 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  14.13 4.32 13.57 4.32 13.57 3.18 12.59 3.18 12.59 2.86
                 13.57 2.86 13.57 1.22 13.89 1.22 13.89 4.00 14.13 4.00 ;
        POLYGON  13.25 2.47 12.93 2.47 12.93 2.28 11.03 2.28 11.03 4.54
                 10.71 4.54 10.71 2.28 10.27 1.84 10.27 1.22 10.59 1.22
                 10.59 1.70 10.85 1.96 13.25 1.96 ;
        RECT  11.49 3.96 12.49 4.28 ;
        RECT  11.09 1.22 12.39 1.54 ;
        RECT  7.37 4.22 10.33 4.54 ;
        POLYGON  10.17 3.90 9.33 3.90 9.33 3.58 9.85 3.58 9.85 2.34 9.69 2.18
                 6.66 2.18 6.66 1.86 9.83 1.86 10.17 2.20 ;
        RECT  7.13 1.22 9.77 1.54 ;
        POLYGON  9.53 2.86 9.21 2.86 9.21 2.82 7.09 2.82 7.09 3.90 6.77 3.90
                 6.77 2.82 4.46 2.82 4.46 3.06 4.14 3.06 4.14 2.50 6.02 2.50
                 6.02 1.22 6.40 1.22 6.40 1.54 6.34 1.54 6.34 2.50 9.53 2.50 ;
        RECT  4.41 3.46 5.45 3.78 ;
        POLYGON  5.09 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 5.09 4.22 ;
        RECT  4.00 1.22 5.00 1.54 ;
        POLYGON  4.03 3.90 3.24 3.90 3.24 3.04 0.80 3.04 0.80 2.66 1.12 2.66
                 1.12 2.72 3.30 2.72 3.30 1.22 3.62 1.22 3.62 3.04 3.56 3.04
                 3.56 3.58 4.03 3.58 ;
        RECT  1.82 1.22 2.92 1.54 ;
        RECT  1.82 3.58 2.92 3.90 ;
    END
END dffnq_4

MACRO dffnq_2
    CLASS CORE ;
    FOREIGN dffnq_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.00 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.03 3.46 8.16 3.46 8.16 3.68 7.84 3.68 7.84 3.14 9.03 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.42 2.08 2.30 2.40 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.81 3.38 14.24 3.38 14.24 2.64 14.25 2.64 14.25 1.64
                 14.57 1.64 14.57 3.06 14.81 3.06 ;
        END
    END q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 0.90 15.27 0.90 15.27 1.66 14.95 1.66 14.95 0.90
                 13.19 0.90 13.19 1.14 12.87 1.14 12.87 0.90 5.70 0.90
                 5.70 1.48 5.38 1.48 5.38 0.90 1.32 0.90 1.32 1.34 1.00 1.34
                 1.00 0.90 0.00 0.90 0.00 -0.90 16.00 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 6.66 0.00 6.66 0.00 4.86 5.94 4.86 5.94 3.74 6.26 3.74
                 6.26 4.86 12.93 4.86 12.93 3.96 13.25 3.96 13.25 4.86
                 15.19 4.86 15.19 4.22 15.51 4.22 15.51 4.86 16.00 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  14.13 4.54 13.57 4.54 13.57 3.18 12.59 3.18 12.59 2.86
                 13.57 2.86 13.57 1.22 13.89 1.22 13.89 4.22 14.13 4.22 ;
        POLYGON  13.25 2.47 12.93 2.47 12.93 2.28 11.03 2.28 11.03 4.54
                 10.71 4.54 10.71 2.28 10.27 1.84 10.27 1.22 10.59 1.22
                 10.59 1.70 10.85 1.96 13.25 1.96 ;
        RECT  11.49 3.96 12.49 4.28 ;
        RECT  11.09 1.22 12.39 1.54 ;
        RECT  7.37 4.22 10.33 4.54 ;
        POLYGON  10.17 3.90 9.33 3.90 9.33 3.58 9.85 3.58 9.85 2.34 9.69 2.18
                 6.66 2.18 6.66 1.86 9.83 1.86 10.17 2.20 ;
        RECT  7.13 1.22 9.77 1.54 ;
        POLYGON  9.53 2.86 9.21 2.86 9.21 2.82 7.09 2.82 7.09 3.90 6.77 3.90
                 6.77 2.82 4.46 2.82 4.46 3.06 4.14 3.06 4.14 2.50 6.02 2.50
                 6.02 1.22 6.40 1.22 6.40 1.54 6.34 1.54 6.34 2.50 9.53 2.50 ;
        RECT  4.41 3.46 5.45 3.78 ;
        POLYGON  5.09 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 5.09 4.22 ;
        RECT  4.00 1.22 5.00 1.54 ;
        POLYGON  4.03 3.90 3.24 3.90 3.24 3.04 0.80 3.04 0.80 2.66 1.12 2.66
                 1.12 2.72 3.30 2.72 3.30 1.22 3.62 1.22 3.62 3.04 3.56 3.04
                 3.56 3.58 4.03 3.58 ;
        RECT  1.82 1.22 2.92 1.54 ;
        RECT  1.82 3.58 2.92 3.90 ;
    END
END dffnq_2

MACRO dffnq_1
    CLASS CORE ;
    FOREIGN dffnq_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.00 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.03 3.46 8.16 3.46 8.16 3.68 7.84 3.68 7.84 3.14 9.03 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.42 2.08 2.30 2.40 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.81 4.18 14.49 4.18 14.49 3.90 14.24 3.90 14.24 3.36
                 14.25 3.36 14.25 1.22 14.57 1.22 14.57 3.58 14.81 3.58 ;
        END
    END q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 0.90 15.27 0.90 15.27 1.24 14.95 1.24 14.95 0.90
                 13.19 0.90 13.19 1.14 12.87 1.14 12.87 0.90 5.70 0.90
                 5.70 1.48 5.38 1.48 5.38 0.90 1.32 0.90 1.32 1.34 1.00 1.34
                 1.00 0.90 0.00 0.90 0.00 -0.90 16.00 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.00 6.66 0.00 6.66 0.00 4.86 5.94 4.86 5.94 3.74 6.26 3.74
                 6.26 4.86 12.93 4.86 12.93 3.96 13.25 3.96 13.25 4.86
                 15.19 4.86 15.19 4.16 15.51 4.16 15.51 4.86 16.00 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  14.13 4.54 13.57 4.54 13.57 3.18 12.59 3.18 12.59 2.86
                 13.57 2.86 13.57 1.22 13.89 1.22 13.89 4.22 14.13 4.22 ;
        POLYGON  13.25 2.47 12.93 2.47 12.93 2.28 11.03 2.28 11.03 4.54
                 10.71 4.54 10.71 2.28 10.27 1.84 10.27 1.22 10.59 1.22
                 10.59 1.70 10.85 1.96 13.25 1.96 ;
        RECT  11.49 3.96 12.49 4.28 ;
        RECT  11.09 1.22 12.39 1.54 ;
        RECT  7.37 4.22 10.33 4.54 ;
        POLYGON  10.17 3.90 9.33 3.90 9.33 3.58 9.85 3.58 9.85 2.34 9.69 2.18
                 6.66 2.18 6.66 1.86 9.83 1.86 10.17 2.20 ;
        RECT  7.13 1.22 9.77 1.54 ;
        POLYGON  9.53 2.86 9.21 2.86 9.21 2.82 7.09 2.82 7.09 3.90 6.77 3.90
                 6.77 2.82 4.46 2.82 4.46 3.06 4.14 3.06 4.14 2.50 6.02 2.50
                 6.02 1.22 6.40 1.22 6.40 1.54 6.34 1.54 6.34 2.50 9.53 2.50 ;
        RECT  4.41 3.46 5.45 3.78 ;
        POLYGON  5.09 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 5.09 4.22 ;
        RECT  4.00 1.22 5.00 1.54 ;
        POLYGON  4.03 3.90 3.24 3.90 3.24 3.04 0.80 3.04 0.80 2.66 1.12 2.66
                 1.12 2.72 3.30 2.72 3.30 1.22 3.62 1.22 3.62 3.04 3.56 3.04
                 3.56 3.58 4.03 3.58 ;
        RECT  1.82 1.22 2.92 1.54 ;
        RECT  1.82 3.58 2.92 3.90 ;
    END
END dffnq_1

MACRO dffn_4
    CLASS CORE ;
    FOREIGN dffn_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.56 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.03 3.46 8.16 3.46 8.16 3.68 7.84 3.68 7.84 3.14 9.03 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.42 2.08 2.30 2.40 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.48 3.26 14.57 3.26 14.57 2.94 16.02 2.94 16.02 1.97
                 14.09 1.97 14.09 1.65 16.34 1.65 16.34 2.72 16.48 2.72 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  18.40 4.54 16.66 4.54 16.66 4.22 18.08 4.22 18.08 1.91
                 16.66 1.91 16.66 1.59 18.40 1.59 ;
        END
    END qb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  18.56 0.90 17.68 0.90 17.68 1.24 17.36 1.24 17.36 0.90
                 15.11 0.90 15.11 1.24 14.79 1.24 14.79 0.90 13.03 0.90
                 13.03 1.14 12.71 1.14 12.71 0.90 5.70 0.90 5.70 1.48 5.38 1.48
                 5.38 0.90 1.32 0.90 1.32 1.34 1.00 1.34 1.00 0.90 0.00 0.90
                 0.00 -0.90 18.56 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  18.56 6.66 0.00 6.66 0.00 4.86 5.94 4.86 5.94 3.74 6.26 3.74
                 6.26 4.86 12.93 4.86 12.93 4.26 13.25 4.26 13.25 4.86
                 15.28 4.86 15.28 4.81 15.60 4.81 15.60 4.86 18.56 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  17.68 3.34 17.25 3.34 17.25 3.90 13.41 3.90 13.41 3.18
                 12.59 3.18 12.59 2.86 13.41 2.86 13.41 1.22 13.73 1.22
                 13.73 3.58 16.93 3.58 16.93 3.02 17.36 3.02 17.36 2.35
                 17.68 2.35 ;
        POLYGON  13.09 2.47 12.77 2.47 12.77 2.28 11.03 2.28 11.03 4.54
                 10.71 4.54 10.71 2.28 10.27 1.84 10.27 1.22 10.59 1.22
                 10.59 1.70 10.85 1.96 13.09 1.96 ;
        RECT  11.49 3.96 12.49 4.28 ;
        RECT  11.09 1.22 12.23 1.54 ;
        RECT  7.37 4.22 10.33 4.54 ;
        POLYGON  10.17 3.90 9.33 3.90 9.33 3.58 9.85 3.58 9.85 2.34 9.69 2.18
                 6.66 2.18 6.66 1.86 9.83 1.86 10.17 2.20 ;
        RECT  7.13 1.22 9.77 1.54 ;
        POLYGON  9.53 2.86 9.21 2.86 9.21 2.82 7.09 2.82 7.09 3.90 6.77 3.90
                 6.77 2.82 4.46 2.82 4.46 3.06 4.14 3.06 4.14 2.50 6.02 2.50
                 6.02 1.22 6.40 1.22 6.40 1.54 6.34 1.54 6.34 2.50 9.53 2.50 ;
        RECT  4.41 3.46 5.45 3.78 ;
        POLYGON  5.09 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 5.09 4.22 ;
        RECT  4.00 1.22 5.00 1.54 ;
        POLYGON  4.03 3.90 3.24 3.90 3.24 3.04 0.80 3.04 0.80 2.66 1.12 2.66
                 1.12 2.72 3.30 2.72 3.30 1.22 3.62 1.22 3.62 3.04 3.56 3.04
                 3.56 3.58 4.03 3.58 ;
        RECT  1.82 1.22 2.92 1.54 ;
        RECT  1.82 3.58 2.92 3.90 ;
    END
END dffn_4

MACRO dffn_2
    CLASS CORE ;
    FOREIGN dffn_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.64 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.03 3.46 8.16 3.46 8.16 3.68 7.84 3.68 7.84 3.14 9.03 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.42 2.08 2.30 2.40 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.82 3.38 14.24 3.38 14.24 2.72 14.50 2.72 14.50 1.64
                 14.82 1.64 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.48 4.44 15.90 4.44 15.90 4.12 16.16 4.12 16.16 1.96
                 15.90 1.96 15.90 1.64 16.48 1.64 ;
        END
    END qb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 0.90 15.52 0.90 15.52 1.24 15.20 1.24 15.20 0.90
                 13.19 0.90 13.19 1.14 12.87 1.14 12.87 0.90 5.70 0.90
                 5.70 1.48 5.38 1.48 5.38 0.90 1.32 0.90 1.32 1.34 1.00 1.34
                 1.00 0.90 0.00 0.90 0.00 -0.90 16.64 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 6.66 0.00 6.66 0.00 4.86 5.94 4.86 5.94 3.74 6.26 3.74
                 6.26 4.86 12.93 4.86 12.93 3.96 13.25 3.96 13.25 4.86
                 16.64 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  15.68 2.68 15.46 2.68 15.46 4.54 13.57 4.54 13.57 3.18
                 12.59 3.18 12.59 2.86 13.57 2.86 13.57 1.22 13.89 1.22
                 13.89 4.22 15.14 4.22 15.14 2.36 15.68 2.36 ;
        POLYGON  13.25 2.47 12.93 2.47 12.93 2.28 11.03 2.28 11.03 4.54
                 10.71 4.54 10.71 2.28 10.27 1.84 10.27 1.22 10.59 1.22
                 10.59 1.70 10.85 1.96 13.25 1.96 ;
        RECT  11.49 3.96 12.49 4.28 ;
        RECT  11.09 1.22 12.39 1.54 ;
        RECT  7.37 4.22 10.33 4.54 ;
        POLYGON  10.17 3.90 9.33 3.90 9.33 3.58 9.85 3.58 9.85 2.34 9.69 2.18
                 6.66 2.18 6.66 1.86 9.83 1.86 10.17 2.20 ;
        RECT  7.13 1.22 9.77 1.54 ;
        POLYGON  9.53 2.86 9.21 2.86 9.21 2.82 7.09 2.82 7.09 3.90 6.77 3.90
                 6.77 2.82 4.46 2.82 4.46 3.06 4.14 3.06 4.14 2.50 6.02 2.50
                 6.02 1.22 6.40 1.22 6.40 1.54 6.34 1.54 6.34 2.50 9.53 2.50 ;
        RECT  4.41 3.46 5.45 3.78 ;
        POLYGON  5.09 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 5.09 4.22 ;
        RECT  4.00 1.22 5.00 1.54 ;
        POLYGON  4.03 3.90 3.24 3.90 3.24 3.04 0.80 3.04 0.80 2.66 1.12 2.66
                 1.12 2.72 3.30 2.72 3.30 1.22 3.62 1.22 3.62 3.04 3.56 3.04
                 3.56 3.58 4.03 3.58 ;
        RECT  1.82 1.22 2.92 1.54 ;
        RECT  1.82 3.58 2.92 3.90 ;
    END
END dffn_2

MACRO dffn_1
    CLASS CORE ;
    FOREIGN dffn_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.64 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.03 3.46 8.16 3.46 8.16 3.68 7.84 3.68 7.84 3.14 9.03 3.14 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.42 2.08 2.30 2.40 ;
        END
    END d
    PIN q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.43  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.81 3.68 14.24 3.68 14.24 3.12 14.25 3.12 14.25 1.22
                 14.57 1.22 14.57 3.34 14.81 3.34 ;
        END
    END q
    PIN qb
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.48 4.08 15.98 4.08 15.98 3.76 16.16 3.76 16.16 1.54
                 15.65 1.54 15.65 1.22 16.48 1.22 ;
        END
    END qb
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 0.90 15.27 0.90 15.27 1.24 14.95 1.24 14.95 0.90
                 13.19 0.90 13.19 1.14 12.87 1.14 12.87 0.90 5.70 0.90
                 5.70 1.48 5.38 1.48 5.38 0.90 1.32 0.90 1.32 1.34 1.00 1.34
                 1.00 0.90 0.00 0.90 0.00 -0.90 16.64 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 6.66 0.00 6.66 0.00 4.86 5.94 4.86 5.94 3.74 6.26 3.74
                 6.26 4.86 12.93 4.86 12.93 3.96 13.25 3.96 13.25 4.86
                 16.64 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  15.45 4.54 13.57 4.54 13.57 3.18 12.59 3.18 12.59 2.86
                 13.57 2.86 13.57 1.22 13.89 1.22 13.89 4.22 15.13 4.22
                 15.13 2.46 15.11 2.46 15.11 2.14 15.45 2.14 ;
        POLYGON  13.25 2.47 12.93 2.47 12.93 2.28 11.03 2.28 11.03 4.54
                 10.71 4.54 10.71 2.28 10.27 1.84 10.27 1.22 10.59 1.22
                 10.59 1.70 10.85 1.96 13.25 1.96 ;
        RECT  11.49 3.96 12.49 4.28 ;
        RECT  11.09 1.22 12.39 1.54 ;
        RECT  7.37 4.22 10.33 4.54 ;
        POLYGON  10.17 3.90 9.33 3.90 9.33 3.58 9.85 3.58 9.85 2.34 9.69 2.18
                 6.66 2.18 6.66 1.86 9.83 1.86 10.17 2.20 ;
        RECT  7.13 1.22 9.77 1.54 ;
        POLYGON  9.53 2.86 9.21 2.86 9.21 2.82 7.09 2.82 7.09 3.90 6.77 3.90
                 6.77 2.82 4.46 2.82 4.46 3.06 4.14 3.06 4.14 2.50 6.02 2.50
                 6.02 1.22 6.40 1.22 6.40 1.54 6.34 1.54 6.34 2.50 9.53 2.50 ;
        RECT  4.41 3.46 5.45 3.78 ;
        POLYGON  5.09 4.54 0.16 4.54 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54
                 0.48 4.22 5.09 4.22 ;
        RECT  4.00 1.22 5.00 1.54 ;
        POLYGON  4.03 3.90 3.24 3.90 3.24 3.04 0.80 3.04 0.80 2.66 1.12 2.66
                 1.12 2.72 3.30 2.72 3.30 1.22 3.62 1.22 3.62 3.04 3.56 3.04
                 3.56 3.58 4.03 3.58 ;
        RECT  1.82 1.22 2.92 1.54 ;
        RECT  1.82 3.58 2.92 3.90 ;
    END
END dffn_1

MACRO dc38_4
    CLASS CORE ;
    FOREIGN dc38_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 117.76 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 10.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  91.65 3.00 90.30 3.00 90.30 4.30 62.56 4.30 62.56 4.32
                 62.14 4.32 62.14 4.30 27.33 4.30 27.33 3.00 25.93 3.00
                 25.93 2.68 27.65 2.68 27.65 3.98 54.44 3.98 54.44 2.67
                 54.76 2.67 54.76 3.98 62.14 3.98 62.14 2.68 62.46 2.68
                 62.46 3.98 89.98 3.98 89.98 2.68 91.65 2.68 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.03  LAYER metal1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 10.15  LAYER metal1  ;
        ANTENNAMAXAREACAR 0.10  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  58.40 2.08 58.72 2.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 10.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  58.08 2.66 56.68 2.66 56.68 2.34 57.76 2.34 57.76 2.08
                 58.08 2.08 ;
        END
    END c
    PIN x0
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.84  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.30 1.72 1.76 1.72 1.76 3.80 3.30 3.80 3.30 4.12 0.18 4.12
                 0.18 3.80 1.44 3.80 1.44 1.72 0.18 1.72 0.18 1.40 3.30 1.40 ;
        END
    END x0
    PIN x1
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.84  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  17.22 1.72 15.84 1.72 15.84 3.42 17.22 3.42 17.22 3.74
                 14.10 3.74 14.10 3.42 15.52 3.42 15.52 1.72 14.10 1.72
                 14.10 1.40 17.22 1.40 ;
        END
    END x1
    PIN x2
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.84  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  31.14 1.60 29.28 1.60 29.28 3.34 31.14 3.34 31.14 3.66
                 28.02 3.66 28.02 3.34 28.96 3.34 28.96 1.60 28.02 1.60
                 28.02 1.28 31.14 1.28 ;
        END
    END x2
    PIN x3
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.84  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  45.06 1.94 43.36 1.94 43.36 3.34 44.58 3.34 44.58 3.66
                 41.46 3.66 41.46 3.34 43.04 3.34 43.04 1.94 41.94 1.94
                 41.94 1.62 45.06 1.62 ;
        END
    END x3
    PIN x4
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.84  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  117.42 1.72 116.32 1.72 116.32 3.80 117.42 3.80 117.42 4.12
                 114.30 4.12 114.30 3.80 116.00 3.80 116.00 1.72 114.30 1.72
                 114.30 1.40 117.42 1.40 ;
        END
    END x4
    PIN x5
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.84  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  103.50 1.72 102.24 1.72 102.24 3.42 103.50 3.42 103.50 3.74
                 100.38 3.74 100.38 3.42 101.92 3.42 101.92 1.72 100.38 1.72
                 100.38 1.40 103.50 1.40 ;
        END
    END x5
    PIN x6
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.84  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  89.58 1.72 88.16 1.72 88.16 3.29 89.58 3.29 89.58 3.61
                 86.46 3.61 86.46 3.29 87.84 3.29 87.84 1.72 86.46 1.72
                 86.46 1.40 89.58 1.40 ;
        END
    END x6
    PIN x7
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.84  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  76.14 3.66 73.02 3.66 73.02 3.34 74.40 3.34 74.40 1.84
                 72.54 1.84 72.54 1.52 75.66 1.52 75.66 1.84 74.72 1.84
                 74.72 3.34 76.14 3.34 ;
        END
    END x7
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  117.76 0.90 78.44 0.90 78.44 1.14 78.12 1.14 78.12 0.90
                 77.04 0.90 77.04 1.14 76.72 1.14 76.72 0.90 74.96 0.90
                 74.96 1.14 74.64 1.14 74.64 0.90 73.56 0.90 73.56 1.14
                 73.24 1.14 73.24 0.90 64.52 0.90 64.52 1.14 64.20 1.14
                 64.20 0.90 63.12 0.90 63.12 1.14 62.80 1.14 62.80 0.90
                 61.04 0.90 61.04 1.14 60.72 1.14 60.72 0.90 56.88 0.90
                 56.88 1.14 56.56 1.14 56.56 0.90 54.80 0.90 54.80 1.14
                 54.48 1.14 54.48 0.90 53.40 0.90 53.40 1.14 53.08 1.14
                 53.08 0.90 44.36 0.90 44.36 1.15 44.04 1.15 44.04 0.90
                 42.96 0.90 42.96 1.15 42.64 1.15 42.64 0.90 40.88 0.90
                 40.88 1.14 40.56 1.14 40.56 0.90 39.48 0.90 39.48 1.14
                 39.16 1.14 39.16 0.90 0.00 0.90 0.00 -0.90 117.76 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  117.76 6.66 0.00 6.66 0.00 4.86 5.04 4.86 5.04 4.62 5.36 4.62
                 5.36 4.86 6.44 4.86 6.44 4.62 6.76 4.62 6.76 4.86 7.84 4.86
                 7.84 4.62 8.16 4.62 8.16 4.86 9.24 4.86 9.24 4.62 9.56 4.62
                 9.56 4.86 10.64 4.86 10.64 4.62 10.96 4.62 10.96 4.86
                 12.04 4.86 12.04 4.62 12.36 4.62 12.36 4.86 14.80 4.86
                 14.80 4.62 15.12 4.62 15.12 4.86 16.20 4.86 16.20 4.62
                 16.52 4.62 16.52 4.86 18.96 4.86 18.96 4.62 19.28 4.62
                 19.28 4.86 20.36 4.86 20.36 4.62 20.68 4.62 20.68 4.86
                 21.76 4.86 21.76 4.62 22.08 4.62 22.08 4.86 23.16 4.86
                 23.16 4.62 23.48 4.62 23.48 4.86 24.56 4.86 24.56 4.62
                 24.88 4.62 24.88 4.86 25.96 4.86 25.96 4.62 26.28 4.62
                 26.28 4.86 28.72 4.86 28.72 4.62 29.04 4.62 29.04 4.86
                 30.12 4.86 30.12 4.62 30.44 4.62 30.44 4.86 32.88 4.86
                 32.88 4.62 33.20 4.62 33.20 4.86 34.28 4.86 34.28 4.62
                 34.60 4.62 34.60 4.86 35.68 4.86 35.68 4.62 36.00 4.62
                 36.00 4.86 37.08 4.86 37.08 4.62 37.40 4.62 37.40 4.86
                 38.48 4.86 38.48 4.62 38.80 4.62 38.80 4.86 39.88 4.86
                 39.88 4.62 40.20 4.62 40.20 4.86 42.16 4.86 42.16 4.62
                 42.48 4.62 42.48 4.86 43.56 4.86 43.56 4.62 43.88 4.62
                 43.88 4.86 46.10 4.86 46.10 4.62 46.42 4.62 46.42 4.86
                 47.50 4.86 47.50 4.62 47.82 4.62 47.82 4.86 48.90 4.86
                 48.90 4.62 49.22 4.62 49.22 4.86 50.30 4.86 50.30 4.62
                 50.62 4.62 50.62 4.86 51.70 4.86 51.70 4.62 52.02 4.62
                 52.02 4.86 53.10 4.86 53.10 4.62 53.42 4.62 53.42 4.86
                 54.50 4.86 54.50 4.62 54.82 4.62 54.82 4.86 56.56 4.86
                 56.56 4.62 56.88 4.62 56.88 4.86 58.64 4.86 58.64 4.62
                 58.96 4.62 58.96 4.86 60.72 4.86 60.72 4.62 61.04 4.62
                 61.04 4.86 63.48 4.86 63.48 4.62 63.80 4.62 63.80 4.86
                 64.88 4.86 64.88 4.62 65.20 4.62 65.20 4.86 66.28 4.86
                 66.28 4.62 66.60 4.62 66.60 4.86 67.68 4.86 67.68 4.62
                 68.00 4.62 68.00 4.86 69.08 4.86 69.08 4.62 69.40 4.62
                 69.40 4.86 70.48 4.86 70.48 4.62 70.80 4.62 70.80 4.86
                 73.72 4.86 73.72 4.62 74.04 4.62 74.04 4.86 75.12 4.86
                 75.12 4.62 75.44 4.62 75.44 4.86 77.40 4.86 77.40 4.62
                 77.72 4.62 77.72 4.86 78.80 4.86 78.80 4.62 79.12 4.62
                 79.12 4.86 80.20 4.86 80.20 4.62 80.52 4.62 80.52 4.86
                 81.60 4.86 81.60 4.62 81.92 4.62 81.92 4.86 83.00 4.86
                 83.00 4.62 83.32 4.62 83.32 4.86 84.40 4.86 84.40 4.62
                 84.72 4.62 84.72 4.86 87.16 4.86 87.16 4.62 87.48 4.62
                 87.48 4.86 88.56 4.86 88.56 4.62 88.88 4.62 88.88 4.86
                 91.32 4.86 91.32 4.62 91.64 4.62 91.64 4.86 92.72 4.86
                 92.72 4.62 93.04 4.62 93.04 4.86 94.12 4.86 94.12 4.62
                 94.44 4.62 94.44 4.86 95.52 4.86 95.52 4.62 95.84 4.62
                 95.84 4.86 96.92 4.86 96.92 4.62 97.24 4.62 97.24 4.86
                 98.32 4.86 98.32 4.62 98.64 4.62 98.64 4.86 101.08 4.86
                 101.08 4.62 101.40 4.62 101.40 4.86 102.48 4.86 102.48 4.62
                 102.80 4.62 102.80 4.86 105.24 4.86 105.24 4.62 105.56 4.62
                 105.56 4.86 106.64 4.86 106.64 4.62 106.96 4.62 106.96 4.86
                 108.04 4.86 108.04 4.62 108.36 4.62 108.36 4.86 109.44 4.86
                 109.44 4.62 109.76 4.62 109.76 4.86 110.84 4.86 110.84 4.62
                 111.16 4.62 111.16 4.86 112.24 4.86 112.24 4.62 112.56 4.62
                 112.56 4.86 117.76 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  115.30 2.68 113.94 2.68 113.94 4.18 104.54 4.18 104.54 3.86
                 113.62 3.86 113.62 2.18 110.82 2.18 110.82 1.86 113.62 1.86
                 113.62 1.22 113.94 1.22 113.94 2.34 115.30 2.34 ;
        POLYGON  113.24 1.54 110.50 1.54 110.50 2.18 107.34 2.18 107.34 1.86
                 110.18 1.86 110.18 1.22 113.24 1.22 ;
        RECT  103.86 1.22 109.76 1.54 ;
        RECT  108.65 2.50 109.05 3.00 ;
        RECT  105.25 2.36 105.57 3.00 ;
        POLYGON  101.38 2.52 100.02 2.52 100.02 4.18 90.62 4.18 90.62 3.86
                 99.70 3.86 99.70 2.18 96.90 2.18 96.90 1.86 99.70 1.86
                 99.70 1.22 100.02 1.22 100.02 2.20 101.38 2.20 ;
        POLYGON  99.32 1.54 96.58 1.54 96.58 2.18 93.42 2.18 93.42 1.86
                 96.26 1.86 96.26 1.22 99.32 1.22 ;
        RECT  89.94 1.22 95.84 1.54 ;
        RECT  94.74 2.50 95.14 3.02 ;
        POLYGON  87.46 2.52 86.10 2.52 86.10 3.66 76.70 3.66 76.70 3.34
                 85.78 3.34 85.78 2.18 82.98 2.18 82.98 1.86 86.10 1.86
                 86.10 2.20 87.46 2.20 ;
        POLYGON  85.40 1.54 82.62 1.54 82.62 2.18 79.50 2.18 79.50 1.86
                 82.30 1.86 82.30 1.22 85.40 1.22 ;
        POLYGON  81.92 1.54 79.14 1.54 79.14 1.80 76.02 1.80 76.02 1.48
                 78.82 1.48 78.82 1.22 81.92 1.22 ;
        RECT  80.82 2.50 81.22 3.00 ;
        RECT  78.11 2.37 78.43 3.00 ;
        POLYGON  73.54 2.66 72.18 2.66 72.18 3.66 62.78 3.66 62.78 3.34
                 71.86 3.34 71.86 2.32 69.06 2.32 69.06 2.00 72.18 2.00
                 72.18 2.34 73.54 2.34 ;
        POLYGON  71.48 1.68 68.74 1.68 68.74 2.18 65.58 2.18 65.58 1.86
                 68.42 1.86 68.42 1.36 71.48 1.36 ;
        POLYGON  68.00 1.54 65.22 1.54 65.22 1.78 62.10 1.78 62.10 1.46
                 64.90 1.46 64.90 1.22 68.00 1.22 ;
        RECT  66.90 2.50 67.30 3.00 ;
        POLYGON  61.74 1.90 60.34 1.90 60.34 3.34 61.74 3.34 61.74 3.66
                 60.02 3.66 60.02 1.44 60.34 1.44 60.34 1.58 61.74 1.58 ;
        POLYGON  59.66 3.66 57.94 3.66 57.94 3.34 59.34 3.34 59.34 1.58
                 57.94 1.58 57.94 1.26 59.66 1.26 ;
        POLYGON  57.58 1.80 56.18 1.80 56.18 3.34 57.58 3.34 57.58 3.66
                 55.08 3.66 55.08 3.34 55.86 3.34 55.86 1.48 57.58 1.48 ;
        POLYGON  55.50 1.78 52.38 1.78 52.38 1.54 49.60 1.54 49.60 1.22
                 52.70 1.22 52.70 1.46 55.50 1.46 ;
        POLYGON  54.12 3.66 45.42 3.66 45.42 2.66 44.06 2.66 44.06 2.34
                 45.42 2.34 45.42 1.86 48.54 1.86 48.54 2.18 45.74 2.18
                 45.74 3.34 54.12 3.34 ;
        POLYGON  52.02 2.18 48.86 2.18 48.86 1.54 46.12 1.54 46.12 1.22
                 49.18 1.22 49.18 1.86 52.02 1.86 ;
        RECT  50.22 2.50 50.62 3.00 ;
        POLYGON  41.58 1.78 38.46 1.78 38.46 1.54 35.68 1.54 35.68 1.22
                 38.78 1.22 38.78 1.46 41.58 1.46 ;
        POLYGON  40.90 3.66 31.50 3.66 31.50 2.54 30.14 2.54 30.14 2.20
                 31.50 2.20 31.50 1.22 31.82 1.22 31.82 1.86 34.62 1.86
                 34.62 2.18 31.82 2.18 31.82 3.34 40.90 3.34 ;
        RECT  39.87 2.36 40.19 3.00 ;
        POLYGON  38.10 2.18 34.94 2.18 34.94 1.54 32.20 1.54 32.20 1.22
                 35.26 1.22 35.26 1.86 38.10 1.86 ;
        RECT  36.30 2.50 36.70 3.00 ;
        RECT  21.76 1.22 27.66 1.54 ;
        POLYGON  26.98 4.20 17.58 4.20 17.58 2.52 16.22 2.52 16.22 2.20
                 17.58 2.20 17.58 1.22 17.90 1.22 17.90 1.86 20.70 1.86
                 20.70 2.18 17.90 2.18 17.90 3.88 26.98 3.88 ;
        POLYGON  24.18 2.18 21.02 2.18 21.02 1.54 18.28 1.54 18.28 1.22
                 21.34 1.22 21.34 1.86 24.18 1.86 ;
        RECT  22.38 2.50 22.78 3.00 ;
        RECT  7.84 1.22 13.74 1.54 ;
        POLYGON  13.06 4.18 3.66 4.18 3.66 2.64 2.30 2.64 2.30 2.32 3.66 2.32
                 3.66 1.22 3.98 1.22 3.98 1.86 6.78 1.86 6.78 2.18 3.98 2.18
                 3.98 3.86 13.06 3.86 ;
        RECT  12.03 2.36 12.35 3.00 ;
        POLYGON  10.26 2.18 7.10 2.18 7.10 1.54 4.36 1.54 4.36 1.22 7.42 1.22
                 7.42 1.86 10.26 1.86 ;
        RECT  8.46 2.50 8.86 3.00 ;
        LAYER v1 ;
        RECT  108.73 2.68 109.05 3.00 ;
        RECT  105.25 2.68 105.57 3.00 ;
        RECT  94.82 2.70 95.14 3.02 ;
        RECT  78.11 2.68 78.43 3.00 ;
        RECT  60.02 1.44 60.34 1.76 ;
        RECT  59.34 3.34 59.66 3.66 ;
        RECT  39.87 2.68 40.19 3.00 ;
        RECT  22.46 2.68 22.78 3.00 ;
        RECT  12.03 2.68 12.35 3.00 ;
        RECT  8.54 2.68 8.86 3.00 ;
        LAYER metal2 ;
        POLYGON  109.05 3.68 8.54 3.68 8.54 2.68 8.86 2.68 8.86 3.36 22.46 3.36
                 22.46 2.68 22.78 2.68 22.78 3.36 59.34 3.36 59.34 3.34
                 59.66 3.34 59.66 3.36 94.82 3.36 94.82 2.70 95.14 2.70
                 95.14 3.36 108.73 3.36 108.73 2.68 109.05 2.68 ;
        POLYGON  105.57 3.00 105.25 3.00 105.25 1.76 78.43 1.76 78.43 3.00
                 78.11 3.00 78.11 1.76 40.19 1.76 40.19 3.00 39.87 3.00
                 39.87 1.76 12.35 1.76 12.35 3.00 12.03 3.00 12.03 1.44
                 105.57 1.44 ;
    END
END dc38_4

MACRO dc38_2
    CLASS CORE ;
    FOREIGN dc38_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 72.96 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN x3
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.04  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  26.86 2.04 25.44 2.04 25.44 3.33 26.38 3.33 26.38 3.65
                 24.66 3.65 24.66 3.33 25.12 3.33 25.12 1.72 26.86 1.72 ;
        END
    END x3
    PIN x4
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.04  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  72.80 4.46 70.90 4.46 70.90 4.14 72.48 4.14 72.48 1.66
                 70.90 1.66 70.90 1.34 72.80 1.34 ;
        END
    END x4
    PIN x5
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.04  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  64.48 4.08 62.58 4.08 62.58 3.76 64.16 3.76 64.16 3.04
                 63.98 3.04 63.98 1.66 62.58 1.66 62.58 1.34 64.30 1.34
                 64.30 2.72 64.48 2.72 ;
        END
    END x5
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 5.54  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  57.38 3.02 56.70 3.02 56.70 4.30 40.16 4.30 40.16 4.32
                 39.84 4.32 39.84 4.30 16.10 4.30 16.10 3.02 15.42 3.02
                 15.42 2.70 16.42 2.70 16.42 3.98 32.04 3.98 32.04 2.70
                 32.36 2.70 32.36 3.98 39.74 3.98 39.74 2.67 40.06 2.67
                 40.06 3.98 56.38 3.98 56.38 2.70 57.38 2.70 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 5.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  36.00 2.08 36.32 2.81 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 5.54  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  35.68 2.56 34.18 2.56 34.18 2.24 35.36 2.24 35.36 2.08
                 35.68 2.08 ;
        END
    END c
    PIN x0
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.04  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.90 1.66 0.48 1.66 0.48 4.14 1.90 4.14 1.90 4.46 0.16 4.46
                 0.16 1.34 1.90 1.34 ;
        END
    END x0
    PIN x1
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.04  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.22 1.66 8.80 1.66 8.80 3.76 10.22 3.76 10.22 4.08 8.48 4.08
                 8.48 1.34 10.22 1.34 ;
        END
    END x1
    PIN x2
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.04  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  18.54 1.66 17.12 1.66 17.12 3.33 18.54 3.33 18.54 3.65
                 16.80 3.65 16.80 1.34 18.54 1.34 ;
        END
    END x2
    PIN x6
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.04  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  55.98 3.65 54.26 3.65 54.26 3.33 55.66 3.33 55.66 1.76
                 54.26 1.76 54.26 1.44 55.98 1.44 ;
        END
    END x6
    PIN x7
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.04  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  48.14 3.66 46.42 3.66 46.42 3.34 47.34 3.34 47.34 2.04
                 45.94 2.04 45.94 1.72 47.66 1.72 47.66 2.72 47.84 2.72
                 47.84 3.34 48.14 3.34 ;
        END
    END x7
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  72.96 0.90 49.04 0.90 49.04 1.14 48.72 1.14 48.72 0.90
                 46.96 0.90 46.96 1.14 46.64 1.14 46.64 0.90 40.72 0.90
                 40.72 1.14 40.40 1.14 40.40 0.90 38.64 0.90 38.64 1.14
                 38.32 1.14 38.32 0.90 34.48 0.90 34.48 1.14 34.16 1.14
                 34.16 0.90 32.40 0.90 32.40 1.14 32.08 1.14 32.08 0.90
                 26.16 0.90 26.16 1.14 25.84 1.14 25.84 0.90 24.08 0.90
                 24.08 1.14 23.76 1.14 23.76 0.90 0.00 0.90 0.00 -0.90
                 72.96 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  72.96 6.66 0.00 6.66 0.00 4.86 3.64 4.86 3.64 4.62 3.96 4.62
                 3.96 4.86 5.04 4.86 5.04 4.62 5.36 4.62 5.36 4.86 6.44 4.86
                 6.44 4.62 6.76 4.62 6.76 4.86 9.20 4.86 9.20 4.62 9.52 4.62
                 9.52 4.86 11.96 4.86 11.96 4.62 12.28 4.62 12.28 4.86
                 13.36 4.86 13.36 4.62 13.68 4.62 13.68 4.86 14.76 4.86
                 14.76 4.62 15.08 4.62 15.08 4.86 17.52 4.86 17.52 4.62
                 17.84 4.62 17.84 4.86 20.28 4.86 20.28 4.62 20.60 4.62
                 20.60 4.86 21.68 4.86 21.68 4.62 22.00 4.62 22.00 4.86
                 23.08 4.86 23.08 4.62 23.40 4.62 23.40 4.86 25.36 4.86
                 25.36 4.62 25.68 4.62 25.68 4.86 27.90 4.86 27.90 4.62
                 28.22 4.62 28.22 4.86 29.30 4.86 29.30 4.62 29.62 4.62
                 29.62 4.86 30.70 4.86 30.70 4.62 31.02 4.62 31.02 4.86
                 32.10 4.86 32.10 4.62 32.42 4.62 32.42 4.86 34.16 4.86
                 34.16 4.62 34.48 4.62 34.48 4.86 36.24 4.86 36.24 4.62
                 36.56 4.62 36.56 4.86 38.32 4.86 38.32 4.62 38.64 4.62
                 38.64 4.86 41.08 4.86 41.08 4.62 41.40 4.62 41.40 4.86
                 42.48 4.86 42.48 4.62 42.80 4.62 42.80 4.86 43.88 4.86
                 43.88 4.62 44.20 4.62 44.20 4.86 47.12 4.86 47.12 4.62
                 47.44 4.62 47.44 4.86 49.40 4.86 49.40 4.62 49.72 4.62
                 49.72 4.86 50.80 4.86 50.80 4.62 51.12 4.62 51.12 4.86
                 52.20 4.86 52.20 4.62 52.52 4.62 52.52 4.86 54.96 4.86
                 54.96 4.62 55.28 4.62 55.28 4.86 57.72 4.86 57.72 4.62
                 58.04 4.62 58.04 4.86 59.12 4.86 59.12 4.62 59.44 4.62
                 59.44 4.86 60.52 4.86 60.52 4.62 60.84 4.62 60.84 4.86
                 63.28 4.86 63.28 4.62 63.60 4.62 63.60 4.86 66.04 4.86
                 66.04 4.62 66.36 4.62 66.36 4.86 67.44 4.86 67.44 4.62
                 67.76 4.62 67.76 4.86 68.84 4.86 68.84 4.62 69.16 4.62
                 69.16 4.86 72.96 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  71.84 2.66 70.54 2.66 70.54 4.18 65.34 4.18 65.34 3.86
                 70.22 3.86 70.22 2.22 68.82 2.22 68.82 1.90 70.54 1.90
                 70.54 2.34 71.84 2.34 ;
        POLYGON  69.84 1.58 68.46 1.58 68.46 2.22 66.74 2.22 66.74 1.90
                 68.14 1.90 68.14 1.26 69.84 1.26 ;
        RECT  64.66 1.26 67.76 1.58 ;
        RECT  67.32 2.54 67.76 3.02 ;
        RECT  65.35 2.38 65.67 3.02 ;
        POLYGON  63.52 2.74 62.22 2.74 62.22 4.18 57.02 4.18 57.02 3.86
                 61.90 3.86 61.90 2.22 60.50 2.22 60.50 1.90 62.22 1.90
                 62.22 2.42 63.52 2.42 ;
        POLYGON  61.52 1.58 60.14 1.58 60.14 2.18 58.42 2.18 58.42 1.86
                 59.82 1.86 59.82 1.26 61.52 1.26 ;
        RECT  56.34 1.22 59.44 1.54 ;
        RECT  58.99 2.54 59.43 3.02 ;
        POLYGON  55.20 2.74 53.90 2.74 53.90 3.66 48.70 3.66 48.70 3.34
                 53.58 3.34 53.58 2.18 52.18 2.18 52.18 1.86 53.90 1.86
                 53.90 2.42 55.20 2.42 ;
        POLYGON  53.20 1.54 51.82 1.54 51.82 2.20 50.10 2.20 50.10 1.88
                 51.50 1.88 51.50 1.22 53.20 1.22 ;
        POLYGON  51.12 1.56 49.74 1.56 49.74 1.90 48.02 1.90 48.02 1.58
                 49.42 1.58 49.42 1.24 51.12 1.24 ;
        RECT  48.72 2.38 49.04 3.02 ;
        POLYGON  46.88 2.68 45.58 2.68 45.58 3.66 40.38 3.66 40.38 3.34
                 45.26 3.34 45.26 2.20 43.86 2.20 43.86 1.88 45.58 1.88
                 45.58 2.36 46.88 2.36 ;
        POLYGON  44.88 1.56 43.50 1.56 43.50 2.20 41.78 2.20 41.78 1.88
                 43.18 1.88 43.18 1.24 44.88 1.24 ;
        POLYGON  42.80 1.56 41.42 1.56 41.42 1.90 39.70 1.90 39.70 1.58
                 41.10 1.58 41.10 1.24 42.80 1.24 ;
        POLYGON  39.34 3.66 37.62 3.66 37.62 3.34 39.02 3.34 39.02 1.90
                 37.62 1.90 37.62 1.58 39.02 1.58 39.02 1.44 39.34 1.44 ;
        POLYGON  37.26 3.66 35.54 3.66 35.54 3.34 36.94 3.34 36.94 1.58
                 35.54 1.58 35.54 1.26 37.26 1.26 ;
        POLYGON  35.18 1.78 33.78 1.78 33.78 3.34 35.18 3.34 35.18 3.66
                 32.68 3.66 32.68 3.34 33.46 3.34 33.46 1.46 35.18 1.46 ;
        POLYGON  33.10 1.90 31.38 1.90 31.38 1.56 30.00 1.56 30.00 1.24
                 31.70 1.24 31.70 1.58 33.10 1.58 ;
        POLYGON  31.72 3.66 27.22 3.66 27.22 2.68 25.92 2.68 25.92 2.36
                 27.22 2.36 27.22 1.88 28.94 1.88 28.94 2.20 27.54 2.20
                 27.54 3.34 31.72 3.34 ;
        POLYGON  31.02 2.20 29.30 2.20 29.30 1.56 27.92 1.56 27.92 1.24
                 29.62 1.24 29.62 1.88 31.02 1.88 ;
        POLYGON  24.78 1.90 23.06 1.90 23.06 1.56 21.68 1.56 21.68 1.24
                 23.38 1.24 23.38 1.58 24.78 1.58 ;
        POLYGON  24.10 3.66 18.90 3.66 18.90 2.74 17.60 2.74 17.60 2.42
                 18.90 2.42 18.90 1.88 20.62 1.88 20.62 2.20 19.22 2.20
                 19.22 3.34 24.10 3.34 ;
        RECT  23.76 2.38 24.08 3.02 ;
        POLYGON  22.70 2.20 20.98 2.20 20.98 1.56 19.60 1.56 19.60 1.24
                 21.30 1.24 21.30 1.88 22.70 1.88 ;
        RECT  13.36 1.22 16.46 1.54 ;
        POLYGON  15.78 4.18 10.58 4.18 10.58 2.74 9.28 2.74 9.28 2.42
                 10.58 2.42 10.58 1.90 12.30 1.90 12.30 2.22 10.90 2.22
                 10.90 3.86 15.78 3.86 ;
        POLYGON  14.38 2.22 12.66 2.22 12.66 1.58 11.28 1.58 11.28 1.26
                 12.98 1.26 12.98 1.90 14.38 1.90 ;
        RECT  13.24 2.54 13.68 3.01 ;
        RECT  5.04 1.26 8.14 1.58 ;
        POLYGON  7.46 4.18 2.26 4.18 2.26 2.66 0.96 2.66 0.96 2.34 2.26 2.34
                 2.26 1.90 3.98 1.90 3.98 2.22 2.58 2.22 2.58 3.86 7.46 3.86 ;
        RECT  7.12 2.38 7.44 3.02 ;
        POLYGON  6.06 2.22 4.34 2.22 4.34 1.58 2.96 1.58 2.96 1.26 4.66 1.26
                 4.66 1.90 6.06 1.90 ;
        RECT  4.92 2.54 5.36 3.02 ;
        LAYER v1 ;
        RECT  67.44 2.70 67.76 3.02 ;
        RECT  65.35 2.70 65.67 3.02 ;
        RECT  59.11 2.70 59.43 3.02 ;
        RECT  48.72 2.70 49.04 3.02 ;
        RECT  39.02 1.44 39.34 1.76 ;
        RECT  36.94 3.34 37.26 3.66 ;
        RECT  23.76 2.70 24.08 3.02 ;
        RECT  13.36 2.69 13.68 3.01 ;
        RECT  7.12 2.70 7.44 3.02 ;
        RECT  5.04 2.70 5.36 3.02 ;
        LAYER metal2 ;
        POLYGON  67.76 3.68 5.04 3.68 5.04 2.70 5.36 2.70 5.36 3.36 13.36 3.36
                 13.36 2.69 13.68 2.69 13.68 3.36 36.94 3.36 36.94 3.34
                 37.26 3.34 37.26 3.36 59.11 3.36 59.11 2.70 59.43 2.70
                 59.43 3.36 67.44 3.36 67.44 2.70 67.76 2.70 ;
        POLYGON  65.67 3.02 65.35 3.02 65.35 1.76 49.04 1.76 49.04 3.02
                 48.72 3.02 48.72 1.76 24.08 1.76 24.08 3.02 23.76 3.02
                 23.76 1.76 7.44 1.76 7.44 3.02 7.12 3.02 7.12 1.44 65.67 1.44 ;
    END
END dc38_2

MACRO dc38_1
    CLASS CORE ;
    FOREIGN dc38_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 44.80 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.79  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  21.24 2.06 21.86 2.40 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.78  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  21.86 3.33 21.54 3.33 21.54 3.04 21.25 3.04 21.25 2.72
                 21.86 2.72 ;
        END
    END c
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.79  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  37.30 4.27 37.29 4.27 37.29 4.30 28.95 4.30 28.95 4.32
                 28.00 4.32 28.00 4.30 22.88 4.30 22.88 4.32 22.56 4.32
                 22.56 4.30 6.60 4.30 6.60 2.78 6.92 2.78 6.92 3.98 16.70 3.98
                 16.70 2.85 17.02 2.85 17.02 3.98 23.50 3.98 23.50 2.90
                 23.83 2.90 23.83 3.98 27.16 3.98 27.16 2.91 26.81 2.91
                 26.81 2.59 27.48 2.59 27.48 3.98 28.17 3.98 28.17 4.00
                 28.79 4.00 28.79 3.98 36.98 3.98 36.98 2.82 37.30 2.82 ;
        END
    END a
    PIN x0
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  0.50 4.11 0.18 4.11 0.18 3.04 0.16 3.04 0.16 2.72 0.18 2.72
                 0.18 1.33 0.50 1.33 ;
        END
    END x0
    PIN x1
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  5.60 3.04 5.58 3.04 5.58 3.83 5.26 3.83 5.26 1.35 5.58 1.35
                 5.58 2.72 5.60 2.72 ;
        END
    END x1
    PIN x2
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.72 3.04 10.66 3.04 10.66 3.48 10.34 3.48 10.34 1.40
                 10.66 1.40 10.66 2.72 10.72 2.72 ;
        END
    END x2
    PIN x3
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  15.74 3.04 15.27 3.04 15.27 3.66 14.88 3.66 14.88 2.72
                 15.42 2.72 15.42 1.66 15.74 1.66 ;
        END
    END x3
    PIN x4
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  44.64 3.04 44.20 3.04 44.20 4.05 43.88 4.05 43.88 1.28
                 44.20 1.28 44.20 2.72 44.64 2.72 ;
        END
    END x4
    PIN x5
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  39.12 4.18 38.32 4.18 38.32 3.86 38.56 3.86 38.56 3.36
                 38.80 3.36 38.80 1.28 39.12 1.28 ;
        END
    END x5
    PIN x6
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  34.04 3.63 33.72 3.63 33.72 1.76 33.44 1.76 33.44 1.27
                 34.04 1.27 ;
        END
    END x6
    PIN x7
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  28.96 3.56 28.64 3.56 28.64 3.68 28.32 3.68 28.32 3.56
                 28.14 3.56 28.14 3.24 28.64 3.24 28.64 1.66 28.96 1.66 ;
        END
    END x7
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  44.80 0.90 28.12 0.90 28.12 1.14 27.80 1.14 27.80 0.90
                 23.88 0.90 23.88 1.22 23.56 1.22 23.56 0.90 21.65 0.90
                 21.65 1.14 21.33 1.14 21.33 0.90 16.58 0.90 16.58 1.14
                 16.26 1.14 16.26 0.90 0.00 0.90 0.00 -0.90 44.80 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  44.80 6.66 0.00 6.66 0.00 4.86 3.88 4.86 3.88 4.62 4.21 4.62
                 4.21 4.86 6.09 4.86 6.09 4.62 6.41 4.62 6.41 4.86 8.96 4.86
                 8.96 4.62 9.29 4.62 9.29 4.86 11.17 4.86 11.17 4.62 11.50 4.62
                 11.50 4.86 13.36 4.86 13.36 4.62 13.69 4.62 13.69 4.86
                 15.77 4.86 15.77 4.62 16.10 4.62 16.10 4.86 18.44 4.86
                 18.44 4.62 18.77 4.62 18.77 4.86 21.48 4.86 21.48 4.62
                 21.80 4.62 21.80 4.86 23.56 4.86 23.56 4.62 23.88 4.62
                 23.88 4.86 24.94 4.86 24.94 4.62 25.26 4.62 25.26 4.86
                 27.32 4.86 27.32 4.62 27.65 4.62 27.65 4.86 30.01 4.86
                 30.01 4.62 30.34 4.62 30.34 4.86 32.88 4.86 32.88 4.62
                 33.21 4.62 33.21 4.86 35.09 4.86 35.09 4.62 35.42 4.62
                 35.42 4.86 37.48 4.86 37.48 4.62 37.81 4.62 37.81 4.86
                 40.17 4.86 40.17 4.62 40.50 4.62 40.50 4.86 44.80 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  43.54 4.28 39.48 4.28 39.48 1.22 39.80 1.22 39.80 3.96
                 43.22 3.96 43.22 2.36 43.54 2.36 ;
        RECT  42.52 2.76 42.84 3.40 ;
        RECT  41.56 1.22 42.56 1.54 ;
        RECT  40.18 1.22 41.18 1.54 ;
        RECT  40.83 2.04 41.15 2.68 ;
        POLYGON  38.44 2.50 36.66 2.50 36.66 3.66 34.40 3.66 34.40 1.24
                 34.72 1.24 34.72 3.34 36.34 3.34 36.34 2.18 38.44 2.18 ;
        RECT  36.48 1.28 37.48 1.60 ;
        RECT  35.10 1.28 36.10 1.60 ;
        RECT  35.70 2.04 36.02 2.68 ;
        POLYGON  33.39 3.66 29.32 3.66 29.32 1.24 29.64 1.24 29.64 3.34
                 33.07 3.34 33.07 2.44 33.39 2.44 ;
        RECT  32.36 2.38 32.68 3.02 ;
        RECT  31.40 1.28 32.40 1.60 ;
        RECT  30.02 1.28 31.02 1.60 ;
        POLYGON  28.32 2.80 28.00 2.80 28.00 2.24 26.49 2.24 26.49 3.34
                 26.84 3.34 26.84 3.66 24.24 3.66 24.24 1.24 24.56 1.24
                 24.56 3.34 26.17 3.34 26.17 1.92 28.32 1.92 ;
        RECT  26.32 1.28 27.32 1.60 ;
        RECT  24.94 1.28 25.94 1.60 ;
        RECT  22.86 1.50 23.18 3.66 ;
        RECT  22.18 1.44 22.50 3.66 ;
        POLYGON  21.10 3.66 20.19 3.66 20.19 3.34 20.46 3.34 20.46 1.58
                 20.83 1.58 20.83 1.90 20.78 1.90 20.78 3.34 21.10 3.34 ;
        POLYGON  20.14 3.01 19.46 3.01 19.46 3.66 17.36 3.66 17.36 2.52
                 16.38 2.52 16.38 2.81 16.06 2.81 16.06 2.20 17.63 2.20
                 17.63 2.25 17.68 2.25 17.68 3.34 19.14 3.34 19.14 2.69
                 19.82 2.69 19.82 1.51 20.14 1.51 ;
        RECT  18.44 1.28 19.44 1.60 ;
        RECT  17.06 1.28 18.06 1.60 ;
        POLYGON  15.06 2.18 14.38 2.18 14.38 3.66 11.12 3.66 11.12 2.44
                 11.44 2.44 11.44 3.34 14.06 3.34 14.06 1.86 14.74 1.86
                 14.74 1.28 15.06 1.28 ;
        RECT  13.36 1.22 14.36 1.54 ;
        RECT  11.98 1.28 12.98 1.60 ;
        RECT  11.76 2.38 12.08 3.02 ;
        POLYGON  9.98 3.66 7.45 3.66 7.45 2.46 6.04 2.46 6.04 2.14 7.77 2.14
                 7.77 3.34 9.66 3.34 9.66 1.28 9.98 1.28 ;
        RECT  8.28 1.28 9.28 1.60 ;
        RECT  8.30 2.04 8.62 2.68 ;
        RECT  6.90 1.28 7.90 1.60 ;
        POLYGON  4.90 4.29 0.95 4.29 0.95 2.36 1.27 2.36 1.27 3.97 4.58 3.97
                 4.58 1.28 4.90 1.28 ;
        RECT  3.20 1.28 4.20 1.60 ;
        RECT  3.17 1.99 3.49 2.66 ;
        RECT  1.82 1.28 2.82 1.60 ;
        RECT  1.59 2.76 1.91 3.40 ;
        LAYER v1 ;
        RECT  42.52 3.08 42.84 3.40 ;
        RECT  40.83 2.36 41.15 2.68 ;
        RECT  35.70 2.36 36.02 2.68 ;
        RECT  32.36 2.70 32.68 3.02 ;
        RECT  22.86 3.34 23.18 3.66 ;
        RECT  22.18 1.44 22.50 1.76 ;
        RECT  11.76 2.70 12.08 3.02 ;
        RECT  8.30 2.36 8.62 2.68 ;
        RECT  3.17 2.34 3.49 2.66 ;
        RECT  1.59 3.08 1.91 3.40 ;
        LAYER metal2 ;
        POLYGON  42.84 3.68 1.59 3.68 1.59 3.08 1.91 3.08 1.91 3.36 11.76 3.36
                 11.76 2.70 12.08 2.70 12.08 3.36 22.86 3.36 22.86 3.34
                 23.18 3.34 23.18 3.36 32.36 3.36 32.36 2.70 32.68 2.70
                 32.68 3.36 42.52 3.36 42.52 3.08 42.84 3.08 ;
        POLYGON  41.15 2.68 40.83 2.68 40.83 1.76 36.02 1.76 36.02 2.68
                 35.70 2.68 35.70 1.76 8.62 1.76 8.62 2.68 8.30 2.68 8.30 1.76
                 3.49 1.76 3.49 2.66 3.17 2.66 3.17 1.44 41.15 1.44 ;
    END
END dc38_1

MACRO dc24_4
    CLASS CORE ;
    FOREIGN dc24_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 47.36 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN x0
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.84  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  46.78 1.74 45.92 1.74 45.92 3.78 46.78 3.78 46.78 4.10
                 43.66 4.10 43.66 3.78 45.60 3.78 45.60 1.74 43.66 1.74
                 43.66 1.42 46.78 1.42 ;
        END
    END x0
    PIN x1
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.84  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.30 1.96 1.90 1.96 1.90 4.00 2.98 4.00 2.98 3.32 3.30 3.32
                 3.30 4.32 0.18 4.32 0.18 3.38 0.50 3.38 0.50 4.00 1.58 4.00
                 1.58 1.96 0.18 1.96 0.18 1.64 3.30 1.64 ;
        END
    END x1
    PIN x2
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.84  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  36.34 1.74 35.04 1.74 35.04 3.58 36.34 3.58 36.34 3.90
                 33.22 3.90 33.22 3.58 34.72 3.58 34.72 1.74 33.22 1.74
                 33.22 1.42 36.34 1.42 ;
        END
    END x2
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 6.54  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  12.44 2.63 13.28 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 6.54  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  22.56 2.62 23.29 3.14 ;
        END
    END b
    PIN x3
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.60  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  15.66 1.78 14.56 1.78 14.56 3.44 15.65 3.44 15.65 3.76
                 13.90 3.76 13.90 3.44 14.24 3.44 14.24 1.78 13.90 1.78
                 13.90 1.46 15.66 1.46 ;
        END
    END x3
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 47.36 6.66 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  47.36 0.90 29.38 0.90 29.38 1.17 29.06 1.17 29.06 0.90
                 27.98 0.90 27.98 1.17 27.66 1.17 27.66 0.90 26.46 0.90
                 26.46 1.19 26.14 1.19 26.14 0.90 24.94 0.90 24.94 1.19
                 24.62 1.19 24.62 0.90 16.34 0.90 16.34 1.14 16.02 1.14
                 16.02 0.90 14.94 0.90 14.94 1.14 14.62 1.14 14.62 0.90
                 13.36 0.90 13.36 1.14 13.04 1.14 13.04 0.90 11.90 0.90
                 11.90 1.14 11.58 1.14 11.58 0.90 10.38 0.90 10.38 1.14
                 10.06 1.14 10.06 0.90 8.86 0.90 8.86 1.14 8.54 1.14 8.54 0.90
                 7.46 0.90 7.46 1.14 7.14 1.14 7.14 0.90 2.60 0.90 2.60 1.18
                 2.28 1.18 2.28 0.90 1.20 0.90 1.20 1.18 0.88 1.18 0.88 0.90
                 0.00 0.90 0.00 -0.90 47.36 -0.90 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        POLYGON  44.60 2.45 43.30 2.45 43.30 4.46 37.38 4.46 37.38 4.14
                 42.98 4.14 42.98 2.22 40.18 2.22 40.18 1.90 42.98 1.90
                 42.98 1.22 43.30 1.22 43.30 2.12 44.60 2.12 ;
        RECT  36.70 1.22 42.60 1.54 ;
        RECT  40.35 2.54 41.17 2.86 ;
        POLYGON  37.80 2.90 37.06 2.90 37.06 4.54 10.23 4.54 10.23 3.26
                 9.27 3.26 9.27 2.94 10.55 2.94 10.55 4.22 25.71 4.22
                 25.71 1.93 23.91 1.93 23.91 1.61 26.03 1.61 26.03 4.22
                 36.74 4.22 36.74 2.58 37.80 2.58 ;
        POLYGON  34.18 2.44 32.86 2.44 32.86 3.90 26.90 3.90 26.90 3.58
                 32.54 3.58 32.54 2.56 29.74 2.56 29.74 2.24 32.54 2.24
                 32.54 1.56 32.86 1.56 32.86 2.12 34.18 2.12 ;
        RECT  26.94 1.49 32.16 1.81 ;
        RECT  28.21 2.13 28.53 3.26 ;
        POLYGON  22.96 3.90 16.70 3.90 16.70 2.66 15.30 2.66 15.30 2.34
                 16.70 2.34 16.70 1.22 17.02 1.22 17.02 1.90 19.82 1.90
                 19.82 2.22 17.02 2.22 17.02 3.58 22.96 3.58 ;
        RECT  17.40 1.22 22.64 1.54 ;
        POLYGON  12.62 1.90 11.90 1.90 11.90 3.58 12.61 3.58 12.61 3.90
                 10.87 3.90 10.87 3.58 11.58 3.58 11.58 1.90 10.87 1.90
                 10.87 1.58 12.62 1.58 ;
        POLYGON  9.83 4.32 3.66 4.32 3.66 2.66 2.37 2.66 2.37 2.34 3.66 2.34
                 3.66 2.16 6.78 2.16 6.78 2.48 3.98 2.48 3.98 4.00 9.83 4.00 ;
        RECT  4.36 1.52 9.58 1.84 ;
        LAYER v1 ;
        RECT  40.85 2.54 41.17 2.86 ;
        RECT  28.21 2.13 28.53 2.45 ;
        RECT  11.58 2.08 11.90 2.40 ;
        LAYER metal2 ;
        POLYGON  41.17 2.86 40.85 2.86 40.85 2.40 28.53 2.40 28.53 2.45
                 28.21 2.45 28.21 2.40 11.58 2.40 11.58 2.08 41.17 2.08 ;
    END
END dc24_4

MACRO dc24_2
    CLASS CORE ;
    FOREIGN dc24_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 27.52 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.27  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  7.32 2.63 8.16 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.27  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  12.64 2.62 13.37 3.14 ;
        END
    END b
    PIN x0
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.04  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  27.36 4.10 25.46 4.10 25.46 3.78 27.04 3.78 27.04 1.74
                 25.46 1.74 25.46 1.42 27.36 1.42 ;
        END
    END x0
    PIN x1
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.04  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.90 1.96 0.50 1.96 0.50 4.00 1.58 4.00 1.58 3.32 1.90 3.32
                 1.90 4.32 0.18 4.32 0.18 1.64 1.90 1.64 ;
        END
    END x1
    PIN x2
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.04  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.96 3.90 19.22 3.90 19.22 3.58 20.62 3.58 20.62 1.74
                 19.22 1.74 19.22 1.42 20.96 1.42 ;
        END
    END x2
    PIN x3
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.80  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.80 3.76 8.32 3.76 8.32 3.44 8.48 3.44 8.48 1.78 8.32 1.78
                 8.32 1.44 8.80 1.44 ;
        END
    END x3
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  27.52 0.90 16.78 0.90 16.78 1.19 16.46 1.19 16.46 0.90
                 15.26 0.90 15.26 1.19 14.94 1.19 14.94 0.90 9.34 0.90
                 9.34 1.14 9.02 1.14 9.02 0.90 7.76 0.90 7.76 1.14 7.44 1.14
                 7.44 0.90 6.26 0.90 6.26 1.14 5.94 1.14 5.94 0.90 4.66 0.90
                 4.66 1.14 4.34 1.14 4.34 0.90 1.20 0.90 1.20 1.18 0.88 1.18
                 0.88 0.90 0.00 0.90 0.00 -0.90 27.52 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 27.52 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  26.40 2.45 25.10 2.45 25.10 4.46 21.97 4.46 21.97 4.14
                 24.78 4.14 24.78 2.22 23.38 2.22 23.38 1.90 25.10 1.90
                 25.10 2.12 26.40 2.12 ;
        RECT  21.30 1.22 24.46 1.54 ;
        RECT  24.05 2.94 24.37 3.68 ;
        POLYGON  22.30 2.90 21.65 2.90 21.65 4.54 6.03 4.54 6.03 3.26 5.07 3.26
                 5.07 2.94 6.35 2.94 6.35 4.22 14.12 4.22 14.12 1.61 14.44 1.61
                 14.44 4.22 21.33 4.22 21.33 2.58 22.30 2.58 ;
        POLYGON  20.18 2.44 18.86 2.44 18.86 3.90 15.69 3.90 15.69 3.58
                 18.50 3.58 18.50 2.56 17.14 2.56 17.14 2.24 18.50 2.24
                 18.50 2.12 20.18 2.12 ;
        RECT  15.75 1.56 18.20 1.88 ;
        POLYGON  15.98 3.26 15.37 3.26 15.37 3.68 15.05 3.68 15.05 2.94
                 15.98 2.94 ;
        POLYGON  13.16 3.90 9.70 3.90 9.70 2.66 9.12 2.66 9.12 2.34 9.70 2.34
                 9.70 1.90 11.42 1.90 11.42 2.22 10.02 2.22 10.02 3.58
                 13.16 3.58 ;
        RECT  10.36 1.22 12.84 1.54 ;
        RECT  6.68 1.58 7.00 3.90 ;
        POLYGON  5.62 4.32 2.29 4.32 2.29 2.66 0.97 2.66 0.97 2.34 2.26 2.34
                 2.26 2.16 3.98 2.16 3.98 2.48 2.61 2.48 2.61 4.00 5.62 4.00 ;
        RECT  2.90 1.52 5.38 1.84 ;
        LAYER v1 ;
        RECT  24.05 3.36 24.37 3.68 ;
        RECT  15.05 3.36 15.37 3.68 ;
        RECT  6.68 3.36 7.00 3.68 ;
        LAYER metal2 ;
        RECT  6.68 3.36 24.37 3.68 ;
    END
END dc24_2

MACRO dc24_1
    CLASS CORE ;
    FOREIGN dc24_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.56 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.26 2.97 3.94 2.97 3.94 2.40 3.36 2.40 3.36 2.08 4.26 2.08 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  8.48 2.08 9.21 2.44 ;
        END
    END b
    PIN x0
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  18.40 4.10 17.97 4.10 17.97 3.78 18.08 3.78 18.08 1.74
                 17.97 1.74 17.97 1.42 18.40 1.42 ;
        END
    END x0
    PIN x1
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 1.64 0.50 4.32 ;
        END
    END x1
    PIN x2
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.15 3.68 13.13 3.68 13.13 3.36 13.83 3.36 13.83 1.42
                 14.15 1.42 ;
        END
    END x2
    PIN x3
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.69  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  5.60 3.68 5.26 3.68 5.26 1.46 5.58 1.46 5.58 3.36 5.60 3.36 ;
        END
    END x3
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  18.56 0.90 11.39 0.90 11.39 1.19 11.07 1.19 11.07 0.90
                 6.28 0.90 6.28 1.14 5.96 1.14 5.96 0.90 4.16 0.90 4.16 1.14
                 3.84 1.14 3.84 0.90 1.20 0.90 1.20 1.18 0.88 1.18 0.88 0.90
                 0.00 0.90 0.00 -0.90 18.56 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 18.56 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  17.76 2.45 16.91 2.45 16.91 4.46 15.21 4.46 15.21 4.14
                 16.59 4.14 16.59 1.59 16.91 1.59 16.91 2.12 17.76 2.12 ;
        RECT  15.18 1.22 16.27 1.54 ;
        RECT  15.82 2.66 16.27 3.26 ;
        POLYGON  14.89 4.54 3.18 4.54 3.18 2.94 3.50 2.94 3.50 4.22 9.65 4.22
                 9.65 1.61 10.00 1.61 10.00 4.22 14.57 4.22 14.57 2.66
                 14.89 2.66 ;
        POLYGON  13.51 2.44 12.77 2.44 12.77 3.90 10.83 3.90 10.83 3.58
                 12.45 3.58 12.45 2.12 13.51 2.12 ;
        RECT  10.36 1.56 12.11 1.88 ;
        RECT  10.53 2.72 11.24 3.04 ;
        POLYGON  8.52 3.90 6.64 3.90 6.64 2.66 5.90 2.66 5.90 2.34 6.64 2.34
                 6.64 1.90 6.96 1.90 6.96 3.58 8.52 3.58 ;
        RECT  7.30 1.22 8.38 1.54 ;
        RECT  4.58 1.57 4.90 3.90 ;
        RECT  2.26 1.43 3.28 1.75 ;
        POLYGON  2.85 4.32 1.56 4.32 1.56 2.66 0.82 2.66 0.82 2.30 1.56 2.30
                 1.56 2.12 1.88 2.12 1.88 4.00 2.85 4.00 ;
        LAYER v1 ;
        RECT  15.95 2.72 16.27 3.04 ;
        RECT  10.92 2.72 11.24 3.04 ;
        RECT  4.58 2.72 4.90 3.04 ;
        LAYER metal2 ;
        RECT  4.58 2.72 16.27 3.04 ;
    END
END dc24_1

MACRO clknor2_8
    CLASS CORE ;
    FOREIGN clknor2_8 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 24.96 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 8.19  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  22.24 2.03 22.97 2.47 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 8.19  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.03 2.00 2.49 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 16.54  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  20.87 1.64 18.07 1.64 18.07 3.21 17.75 3.21 17.75 1.64
                 12.47 1.64 12.47 2.89 17.75 2.89 17.75 3.21 12.15 3.21
                 12.15 1.64 6.91 1.64 6.91 2.89 12.15 2.89 12.15 3.21 6.54 3.21
                 6.54 1.64 3.75 1.64 3.75 1.32 20.87 1.32 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 24.96 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  24.96 6.66 0.00 6.66 0.00 4.85 0.97 4.85 0.97 3.84 1.29 3.84
                 1.29 4.85 2.37 4.85 2.37 3.84 2.69 3.84 2.69 4.85 3.77 4.85
                 3.77 3.86 4.09 3.86 4.09 4.85 5.17 4.85 5.17 3.86 5.49 3.86
                 5.49 4.85 19.13 4.85 19.13 4.51 19.45 4.51 19.45 4.85
                 20.53 4.85 20.53 4.51 20.85 4.51 20.85 4.85 21.93 4.85
                 21.93 4.49 22.25 4.49 22.25 4.85 23.33 4.85 23.33 4.49
                 23.65 4.49 23.65 4.85 24.96 4.85 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  24.35 4.14 18.75 4.14 18.75 4.53 7.19 4.53 7.19 4.21
                 18.43 4.21 18.43 3.13 18.75 3.13 18.75 3.82 19.82 3.82
                 19.82 3.12 20.16 3.12 20.16 3.82 21.22 3.82 21.22 3.12
                 21.56 3.12 21.56 3.82 22.63 3.82 22.63 3.13 22.95 3.13
                 22.95 3.82 24.03 3.82 24.03 3.13 24.35 3.13 ;
        POLYGON  17.40 3.85 5.87 3.85 5.87 3.37 4.79 3.37 4.79 4.20 4.47 4.20
                 4.47 3.37 3.39 3.37 3.39 4.20 3.07 4.20 3.07 3.37 1.99 3.37
                 1.99 4.19 1.67 4.19 1.67 3.37 0.59 3.37 0.59 4.19 0.27 4.19
                 0.27 3.05 6.19 3.05 6.19 3.53 17.40 3.53 ;
    END
END clknor2_8

MACRO clknor2_4
    CLASS CORE ;
    FOREIGN clknor2_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 13.44 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 4.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  11.04 2.04 11.77 2.48 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 4.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.04 2.00 2.57 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 8.83  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  11.06 1.69 9.66 1.69 9.66 3.22 9.34 3.22 9.34 1.69 6.88 1.69
                 6.88 2.90 9.34 2.90 9.34 3.22 6.56 3.22 6.56 1.69 4.06 1.69
                 4.06 2.90 6.56 2.90 6.56 3.22 3.74 3.22 3.74 1.69 2.33 1.69
                 2.33 1.37 11.06 1.37 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 13.44 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  13.44 6.66 0.00 6.66 0.00 4.86 0.96 4.86 0.96 3.85 1.28 3.85
                 1.28 4.86 2.36 4.86 2.36 3.85 2.68 3.85 2.68 4.86 10.72 4.86
                 10.72 4.50 11.04 4.50 11.04 4.86 12.12 4.86 12.12 4.50
                 12.44 4.50 12.44 4.86 13.44 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  13.14 4.15 10.34 4.15 10.34 4.54 4.34 4.54 4.34 4.22
                 10.02 4.22 10.02 3.14 10.34 3.14 10.34 3.83 11.42 3.83
                 11.42 3.14 11.74 3.14 11.74 3.83 12.82 3.83 12.82 3.14
                 13.14 3.14 ;
        POLYGON  8.99 3.86 3.06 3.86 3.06 3.38 1.98 3.38 1.98 4.20 1.66 4.20
                 1.66 3.38 0.58 3.38 0.58 4.20 0.26 4.20 0.26 3.06 3.38 3.06
                 3.38 3.54 8.99 3.54 ;
    END
END clknor2_4

MACRO clknor2_2
    CLASS CORE ;
    FOREIGN clknor2_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.05  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.23 2.04 6.94 2.48 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.05  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.75 2.04 1.29 2.57 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  5.39 1.69 4.32 1.69 4.32 2.90 5.39 2.90 5.39 3.22 2.26 3.22
                 2.26 2.90 4.00 2.90 4.00 1.69 2.26 1.69 2.26 1.37 5.39 1.37 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 7.68 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 7.68 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  7.46 4.49 7.14 4.49 7.14 3.80 6.06 3.80 6.06 4.54 2.94 4.54
                 2.94 4.22 5.74 4.22 5.74 3.48 7.46 3.48 ;
        POLYGON  4.70 3.86 1.58 3.86 1.58 3.72 0.50 3.72 0.50 4.54 0.18 4.54
                 0.18 3.40 1.90 3.40 1.90 3.54 4.70 3.54 ;
    END
END clknor2_2

MACRO clknor2_1
    CLASS CORE ;
    FOREIGN clknor2_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.96  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.08 4.05 2.52 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.96  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.42 2.61 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.75  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  2.69 3.22 2.37 3.22 2.37 1.88 2.08 1.88 2.08 1.42 2.69 1.42 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 5.12 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 6.66 0.00 6.66 0.00 4.86 0.99 4.86 0.99 3.85 1.31 3.85
                 1.31 4.86 5.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.85 4.15 4.22 4.15 4.22 4.54 1.67 4.54 1.67 4.22 3.90 4.22
                 3.90 3.83 4.53 3.83 4.53 3.14 4.85 3.14 ;
        POLYGON  3.43 3.86 1.69 3.86 1.69 3.38 0.61 3.38 0.61 4.20 0.29 4.20
                 0.29 3.06 2.01 3.06 2.01 3.54 3.43 3.54 ;
    END
END clknor2_1

MACRO clknand2_8
    CLASS CORE ;
    FOREIGN clknand2_8 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 24.96 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 8.01  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.49 2.62 7.12 3.19 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 8.01  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  14.24 3.10 14.81 3.69 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 18.47  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  23.24 4.54 12.32 4.54 12.32 2.22 9.57 2.22 9.57 4.22
                 12.32 4.22 12.32 4.54 0.46 4.54 0.46 4.22 9.25 4.22 9.25 2.22
                 6.46 2.22 6.46 1.90 17.98 1.90 17.98 2.22 12.64 2.22
                 12.64 4.22 23.24 4.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 24.96 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 24.96 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  12.75 1.22 24.27 1.54 ;
        RECT  0.18 1.22 11.68 1.54 ;
    END
END clknand2_8

MACRO clknand2_4
    CLASS CORE ;
    FOREIGN clknand2_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 13.44 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 4.00  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 2.62 5.91 3.19 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 4.00  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  8.87 3.10 9.44 3.69 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 9.70  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.04 4.54 7.20 4.54 7.20 2.22 3.97 2.22 3.97 4.22 7.20 4.22
                 7.20 4.54 0.52 4.54 0.52 4.22 3.65 4.22 3.65 1.90 9.59 1.90
                 9.59 2.22 7.52 2.22 7.52 4.22 12.04 4.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 13.44 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 13.44 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  7.15 1.22 13.06 1.54 ;
        RECT  0.18 1.22 6.08 1.54 ;
    END
END clknand2_4

MACRO clknand2_2
    CLASS CORE ;
    FOREIGN clknand2_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.00  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.48 2.62 3.11 3.19 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.00  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.83 3.10 6.40 3.69 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.35  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  6.44 4.54 4.64 4.54 4.64 2.22 1.17 2.22 1.17 4.22 4.64 4.22
                 4.64 4.54 0.52 4.54 0.52 4.22 0.85 4.22 0.85 1.90 5.38 1.90
                 5.38 2.22 4.96 2.22 4.96 4.22 6.44 4.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 7.68 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 7.68 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  4.35 1.22 7.46 1.54 ;
        RECT  0.17 1.22 3.28 1.54 ;
    END
END clknand2_2

MACRO clknand2_1
    CLASS CORE ;
    FOREIGN clknand2_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.00  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.39 2.62 2.02 3.19 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.00  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.99 3.27 3.68 3.75 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.32 4.54 0.85 4.54 0.85 4.22 4.00 4.22 4.00 2.22 2.25 2.22
                 2.25 1.90 4.32 1.90 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 0.90 3.97 0.90 3.97 0.94 3.63 0.94 3.63 0.90 1.21 0.90
                 1.21 0.94 0.87 0.94 0.87 0.90 0.00 0.90 0.00 -0.90 5.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 5.12 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  2.96 1.26 4.66 1.58 ;
        RECT  0.17 1.26 1.88 1.58 ;
    END
END clknand2_1

MACRO clkmux2_4
    CLASS CORE ;
    FOREIGN clkmux2_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.72 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  9.76 2.50 10.08 3.20 ;
        END
    END d0
    PIN d1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.78 ;
        END
    END d1
    PIN sl0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.34  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 1.92 5.60 2.62 ;
        END
    END sl0
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.55  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.56 4.54 14.15 4.54 14.15 3.98 13.07 3.98 13.07 4.54
                 12.75 4.54 12.75 3.98 11.67 3.98 11.67 4.54 11.35 4.54
                 11.35 3.66 14.24 3.66 14.24 1.54 11.35 1.54 11.35 1.22
                 14.56 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 14.72 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  14.72 6.66 0.00 6.66 0.00 4.86 12.05 4.86 12.05 4.30
                 12.37 4.30 12.37 4.86 13.45 4.86 13.45 4.30 13.77 4.30
                 13.77 4.86 14.72 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  12.98 2.69 11.01 2.69 11.01 2.18 8.91 2.18 8.91 3.26 7.03 3.26
                 7.03 2.94 8.59 2.94 8.59 2.18 7.11 2.18 7.11 1.54 4.14 1.54
                 4.14 3.26 3.82 3.26 3.82 2.18 2.58 2.18 2.58 3.26 2.26 3.26
                 2.26 1.86 3.82 1.86 3.82 1.22 7.43 1.22 7.43 1.86 11.33 1.86
                 11.33 2.36 12.98 2.36 ;
        RECT  7.80 1.22 11.02 1.54 ;
        RECT  3.01 3.58 10.99 3.90 ;
        RECT  0.18 4.22 8.18 4.54 ;
        POLYGON  6.78 2.72 6.38 2.72 6.38 3.26 4.50 3.26 4.50 1.86 4.82 1.86
                 4.82 2.94 6.06 2.94 6.06 1.86 6.38 1.86 6.38 2.40 6.78 2.40 ;
        RECT  0.18 1.22 3.37 1.54 ;
    END
END clkmux2_4

MACRO clkmux2_2
    CLASS CORE ;
    FOREIGN clkmux2_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.96 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 1.96 5.60 2.60 ;
        END
    END d0
    PIN d1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.92 1.96 6.24 2.60 ;
        END
    END d1
    PIN sl0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.17  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.72 1.44 3.04 ;
        END
    END sl0
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.86  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.65 4.54 8.33 4.54 8.33 3.98 7.25 3.98 7.25 4.54 6.93 4.54
                 6.93 3.66 8.33 3.66 8.33 2.40 7.84 2.40 7.84 2.08 8.33 2.08
                 8.33 1.54 6.93 1.54 6.93 1.22 8.65 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.96 0.90 1.20 0.90 1.20 1.00 0.88 1.00 0.88 0.90 0.00 0.90
                 0.00 -0.90 8.96 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  8.96 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 5.34 4.86 5.34 4.22 5.66 4.22 5.66 4.86 7.63 4.86
                 7.63 4.30 7.95 4.30 7.95 4.86 8.96 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  7.31 3.24 3.38 3.24 3.38 3.42 3.06 3.42 3.06 2.18 2.39 2.18
                 2.39 1.86 3.38 1.86 3.38 2.92 7.31 2.92 ;
        RECT  1.56 1.22 6.57 1.54 ;
        POLYGON  6.57 4.54 6.25 4.54 6.25 3.90 3.76 3.90 3.76 3.58 6.57 3.58 ;
        RECT  3.76 1.86 4.96 2.18 ;
        RECT  1.56 4.22 4.76 4.54 ;
        POLYGON  2.74 3.90 0.50 3.90 0.50 4.06 0.16 4.06 0.16 1.44 0.50 1.44
                 0.50 1.76 0.48 1.76 0.48 3.58 2.42 3.58 2.42 2.62 2.74 2.62 ;
    END
END clkmux2_2

MACRO clkmux2_1
    CLASS CORE ;
    FOREIGN clkmux2_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.32 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN d0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 1.98 5.60 2.62 ;
        END
    END d0
    PIN d1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.92 1.98 6.24 2.62 ;
        END
    END d1
    PIN sl0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.17  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.72 1.44 3.04 ;
        END
    END sl0
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.43  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.16 2.40 7.95 2.40 7.95 3.72 7.63 3.72 7.63 1.41 7.95 1.41
                 7.95 2.08 8.16 2.08 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 0.90 1.20 0.90 1.20 1.00 0.88 1.00 0.88 0.90 0.00 0.90
                 0.00 -0.90 8.32 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 5.34 4.86 5.34 4.22 5.66 4.22 5.66 4.86 6.93 4.86
                 6.93 4.14 7.25 4.14 7.25 4.86 8.32 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  7.31 3.26 3.38 3.26 3.38 3.42 3.06 3.42 3.06 2.18 2.39 2.18
                 2.39 1.86 3.38 1.86 3.38 2.94 6.99 2.94 6.99 2.59 7.31 2.59 ;
        RECT  1.56 1.22 6.57 1.54 ;
        POLYGON  6.57 4.46 6.25 4.46 6.25 3.90 3.76 3.90 3.76 3.58 6.57 3.58 ;
        RECT  3.76 1.86 4.96 2.18 ;
        RECT  1.56 4.22 4.76 4.54 ;
        POLYGON  2.74 3.90 0.50 3.90 0.50 4.06 0.16 4.06 0.16 1.44 0.50 1.44
                 0.50 1.76 0.48 1.76 0.48 3.58 2.42 3.58 2.42 2.62 2.74 2.62 ;
    END
END clkmux2_1

MACRO clkinv_8
    CLASS CORE ;
    FOREIGN clkinv_8 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 4.98  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.34 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 8.44  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  6.10 1.96 4.70 1.96 4.70 2.72 4.96 2.72 4.96 3.04 4.70 3.04
                 4.70 3.78 6.10 3.78 6.10 4.10 4.38 4.10 4.38 1.96 1.90 1.96
                 1.90 3.78 4.38 3.78 4.38 4.10 0.18 4.10 0.18 3.78 1.58 3.78
                 1.58 1.96 0.18 1.96 0.18 1.64 6.10 1.64 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 0.90 5.40 0.90 5.40 1.32 5.08 1.32 5.08 0.90 4.00 0.90
                 4.00 1.32 3.68 1.32 3.68 0.90 2.60 0.90 2.60 1.32 2.28 1.32
                 2.28 0.90 1.20 0.90 1.20 1.32 0.88 1.32 0.88 0.90 0.00 0.90
                 0.00 -0.90 6.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.42 1.20 4.42
                 1.20 4.86 2.28 4.86 2.28 4.42 2.60 4.42 2.60 4.86 3.68 4.86
                 3.68 4.42 4.00 4.42 4.00 4.86 5.08 4.86 5.08 4.42 5.40 4.42
                 5.40 4.86 6.40 4.86 ;
        END
    END vdd!
END clkinv_8

MACRO clkinv_64
    CLASS CORE ;
    FOREIGN clkinv_64 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 46.08 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 39.86  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.34 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 58.82  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  45.30 1.96 43.90 1.96 43.90 2.72 44.00 2.72 44.00 3.22
                 43.90 3.22 43.90 3.96 44.98 3.96 44.98 3.34 45.30 3.34
                 45.30 4.28 43.58 4.28 43.58 1.96 41.10 1.96 41.10 3.96
                 42.18 3.96 42.18 3.28 42.50 3.28 42.50 3.96 43.58 3.96
                 43.58 4.28 40.78 4.28 40.78 1.96 38.30 1.96 38.30 3.96
                 39.38 3.96 39.38 3.34 39.70 3.34 39.70 3.96 40.78 3.96
                 40.78 4.28 37.98 4.28 37.98 1.96 35.50 1.96 35.50 3.96
                 36.58 3.96 36.58 3.28 36.90 3.28 36.90 3.96 37.98 3.96
                 37.98 4.28 35.18 4.28 35.18 1.96 32.70 1.96 32.70 3.96
                 33.78 3.96 33.78 3.34 34.10 3.34 34.10 3.96 35.18 3.96
                 35.18 4.28 32.38 4.28 32.38 1.96 29.90 1.96 29.90 3.96
                 30.98 3.96 30.98 3.28 31.30 3.28 31.30 3.96 32.38 3.96
                 32.38 4.28 29.58 4.28 29.58 1.96 27.10 1.96 27.10 3.96
                 28.18 3.96 28.18 3.34 28.50 3.34 28.50 3.96 29.58 3.96
                 29.58 4.28 26.78 4.28 26.78 1.96 24.30 1.96 24.30 3.96
                 25.38 3.96 25.38 3.28 25.70 3.28 25.70 3.96 26.78 3.96
                 26.78 4.28 23.98 4.28 23.98 1.96 21.50 1.96 21.50 3.96
                 22.58 3.96 22.58 3.34 22.90 3.34 22.90 3.96 23.98 3.96
                 23.98 4.28 21.18 4.28 21.18 1.96 18.70 1.96 18.70 3.96
                 19.78 3.96 19.78 3.28 20.10 3.28 20.10 3.96 21.18 3.96
                 21.18 4.28 18.38 4.28 18.38 1.96 15.90 1.96 15.90 3.96
                 16.98 3.96 16.98 3.34 17.30 3.34 17.30 3.96 18.38 3.96
                 18.38 4.28 15.58 4.28 15.58 1.96 13.10 1.96 13.10 3.96
                 14.18 3.96 14.18 3.28 14.50 3.28 14.50 3.96 15.58 3.96
                 15.58 4.28 12.78 4.28 12.78 1.96 10.30 1.96 10.30 3.96
                 11.38 3.96 11.38 3.34 11.70 3.34 11.70 3.96 12.78 3.96
                 12.78 4.28 9.98 4.28 9.98 1.96 7.50 1.96 7.50 3.96 8.58 3.96
                 8.58 3.28 8.90 3.28 8.90 3.96 9.98 3.96 9.98 4.28 7.18 4.28
                 7.18 1.96 4.70 1.96 4.70 3.96 5.78 3.96 5.78 3.34 6.10 3.34
                 6.10 3.96 7.18 3.96 7.18 4.28 4.38 4.28 4.38 1.96 1.90 1.96
                 1.90 3.96 2.98 3.96 2.98 3.28 3.30 3.28 3.30 3.96 4.38 3.96
                 4.38 4.28 0.18 4.28 0.18 3.34 0.50 3.34 0.50 3.96 1.58 3.96
                 1.58 1.96 0.18 1.96 0.18 1.64 45.30 1.64 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  46.08 0.90 44.60 0.90 44.60 1.32 44.28 1.32 44.28 0.90
                 43.20 0.90 43.20 1.32 42.88 1.32 42.88 0.90 41.80 0.90
                 41.80 1.32 41.48 1.32 41.48 0.90 40.40 0.90 40.40 1.32
                 40.08 1.32 40.08 0.90 39.00 0.90 39.00 1.32 38.68 1.32
                 38.68 0.90 37.60 0.90 37.60 1.32 37.28 1.32 37.28 0.90
                 36.20 0.90 36.20 1.32 35.88 1.32 35.88 0.90 34.80 0.90
                 34.80 1.32 34.48 1.32 34.48 0.90 33.40 0.90 33.40 1.32
                 33.08 1.32 33.08 0.90 32.00 0.90 32.00 1.32 31.68 1.32
                 31.68 0.90 30.60 0.90 30.60 1.32 30.28 1.32 30.28 0.90
                 29.20 0.90 29.20 1.32 28.88 1.32 28.88 0.90 27.80 0.90
                 27.80 1.32 27.48 1.32 27.48 0.90 26.40 0.90 26.40 1.32
                 26.08 1.32 26.08 0.90 25.00 0.90 25.00 1.32 24.68 1.32
                 24.68 0.90 23.60 0.90 23.60 1.32 23.28 1.32 23.28 0.90
                 22.20 0.90 22.20 1.32 21.88 1.32 21.88 0.90 20.80 0.90
                 20.80 1.32 20.48 1.32 20.48 0.90 19.40 0.90 19.40 1.32
                 19.08 1.32 19.08 0.90 18.00 0.90 18.00 1.32 17.68 1.32
                 17.68 0.90 16.60 0.90 16.60 1.32 16.28 1.32 16.28 0.90
                 15.20 0.90 15.20 1.32 14.88 1.32 14.88 0.90 13.80 0.90
                 13.80 1.32 13.48 1.32 13.48 0.90 12.40 0.90 12.40 1.32
                 12.08 1.32 12.08 0.90 11.00 0.90 11.00 1.32 10.68 1.32
                 10.68 0.90 9.60 0.90 9.60 1.32 9.28 1.32 9.28 0.90 8.20 0.90
                 8.20 1.32 7.88 1.32 7.88 0.90 6.80 0.90 6.80 1.32 6.48 1.32
                 6.48 0.90 5.40 0.90 5.40 1.32 5.08 1.32 5.08 0.90 4.00 0.90
                 4.00 1.32 3.68 1.32 3.68 0.90 2.60 0.90 2.60 1.32 2.28 1.32
                 2.28 0.90 1.20 0.90 1.20 1.32 0.88 1.32 0.88 0.90 0.00 0.90
                 0.00 -0.90 46.08 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 46.08 6.66 ;
        END
    END vdd!
END clkinv_64

MACRO clkinv_6
    CLASS CORE ;
    FOREIGN clkinv_6 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.64  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.70 1.96 3.30 1.96 3.30 3.56 4.38 3.56 4.38 3.34 4.70 3.34
                 4.70 4.38 4.38 4.38 4.38 3.88 3.30 3.88 3.30 4.38 2.98 4.38
                 2.98 3.04 2.72 3.04 2.72 2.72 2.98 2.72 2.98 1.96 1.90 1.96
                 1.90 3.56 2.98 3.56 2.98 3.88 1.90 3.88 1.90 4.38 1.58 4.38
                 1.58 3.88 0.50 3.88 0.50 4.38 0.18 4.38 0.18 3.34 0.50 3.34
                 0.50 3.56 1.58 3.56 1.58 1.96 0.18 1.96 0.18 1.64 4.70 1.64 ;
        END
    END x
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.74  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.34 1.12 3.04 ;
        END
    END a
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.34 1.20 4.34
                 1.20 4.86 2.28 4.86 2.28 4.34 2.60 4.34 2.60 4.86 3.68 4.86
                 3.68 4.34 4.00 4.34 4.00 4.86 5.12 4.86 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 0.90 4.00 0.90 4.00 1.32 3.68 1.32 3.68 0.90 2.60 0.90
                 2.60 1.32 2.28 1.32 2.28 0.90 1.20 0.90 1.20 1.32 0.88 1.32
                 0.88 0.90 0.00 0.90 0.00 -0.90 5.12 -0.90 ;
        END
    END gnd!
END clkinv_6

MACRO clkinv_48
    CLASS CORE ;
    FOREIGN clkinv_48 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 34.56 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 29.89  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.34 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 44.43  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  34.10 1.96 32.70 1.96 32.70 3.56 33.78 3.56 33.78 3.34
                 34.10 3.34 34.10 4.38 33.78 4.38 33.78 3.88 32.70 3.88
                 32.70 4.38 32.38 4.38 32.38 3.11 32.16 3.11 32.16 2.72
                 32.38 2.72 32.38 1.96 31.30 1.96 31.30 3.56 32.38 3.56
                 32.38 3.88 31.30 3.88 31.30 4.38 30.98 4.38 30.98 1.96
                 28.50 1.96 28.50 3.56 29.58 3.56 29.58 3.34 29.90 3.34
                 29.90 3.56 30.98 3.56 30.98 3.88 29.90 3.88 29.90 4.38
                 29.58 4.38 29.58 3.88 28.50 3.88 28.50 4.38 28.18 4.38
                 28.18 1.96 27.10 1.96 27.10 3.56 28.18 3.56 28.18 3.88
                 27.10 3.88 27.10 4.38 26.78 4.38 26.78 1.96 24.30 1.96
                 24.30 3.56 25.38 3.56 25.38 3.34 25.70 3.34 25.70 3.56
                 26.78 3.56 26.78 3.88 25.70 3.88 25.70 4.38 25.38 4.38
                 25.38 3.88 24.30 3.88 24.30 4.38 23.98 4.38 23.98 1.96
                 22.90 1.96 22.90 3.56 23.98 3.56 23.98 3.88 22.90 3.88
                 22.90 4.38 22.58 4.38 22.58 1.96 20.10 1.96 20.10 3.56
                 21.18 3.56 21.18 3.34 21.50 3.34 21.50 3.56 22.58 3.56
                 22.58 3.88 21.50 3.88 21.50 4.38 21.18 4.38 21.18 3.88
                 20.10 3.88 20.10 4.38 19.78 4.38 19.78 1.96 18.70 1.96
                 18.70 3.56 19.78 3.56 19.78 3.88 18.70 3.88 18.70 4.38
                 18.38 4.38 18.38 1.96 15.90 1.96 15.90 3.56 16.98 3.56
                 16.98 3.34 17.30 3.34 17.30 3.56 18.38 3.56 18.38 3.88
                 17.30 3.88 17.30 4.38 16.98 4.38 16.98 3.88 15.90 3.88
                 15.90 4.38 15.58 4.38 15.58 1.96 14.50 1.96 14.50 3.56
                 15.58 3.56 15.58 3.88 14.50 3.88 14.50 4.38 14.18 4.38
                 14.18 1.96 11.70 1.96 11.70 3.56 12.78 3.56 12.78 3.34
                 13.10 3.34 13.10 3.56 14.18 3.56 14.18 3.88 13.10 3.88
                 13.10 4.38 12.78 4.38 12.78 3.88 11.70 3.88 11.70 4.38
                 11.38 4.38 11.38 1.96 10.30 1.96 10.30 3.56 11.38 3.56
                 11.38 3.88 10.30 3.88 10.30 4.38 9.98 4.38 9.98 1.96 7.50 1.96
                 7.50 3.56 8.58 3.56 8.58 3.34 8.90 3.34 8.90 3.56 9.98 3.56
                 9.98 3.88 8.90 3.88 8.90 4.38 8.58 4.38 8.58 3.88 7.50 3.88
                 7.50 4.38 7.18 4.38 7.18 1.96 6.10 1.96 6.10 3.56 7.18 3.56
                 7.18 3.88 6.10 3.88 6.10 4.38 5.78 4.38 5.78 1.96 3.30 1.96
                 3.30 3.56 4.38 3.56 4.38 3.34 4.70 3.34 4.70 3.56 5.78 3.56
                 5.78 3.88 4.70 3.88 4.70 4.38 4.38 4.38 4.38 3.88 3.30 3.88
                 3.30 4.38 2.98 4.38 2.98 1.96 1.90 1.96 1.90 3.56 2.98 3.56
                 2.98 3.88 1.90 3.88 1.90 4.38 1.58 4.38 1.58 3.88 0.50 3.88
                 0.50 4.38 0.18 4.38 0.18 3.34 0.50 3.34 0.50 3.56 1.58 3.56
                 1.58 1.96 0.18 1.96 0.18 1.64 34.10 1.64 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  34.56 0.90 33.40 0.90 33.40 1.32 33.08 1.32 33.08 0.90
                 32.00 0.90 32.00 1.32 31.68 1.32 31.68 0.90 30.60 0.90
                 30.60 1.32 30.28 1.32 30.28 0.90 29.20 0.90 29.20 1.32
                 28.88 1.32 28.88 0.90 27.80 0.90 27.80 1.32 27.48 1.32
                 27.48 0.90 26.40 0.90 26.40 1.32 26.08 1.32 26.08 0.90
                 25.00 0.90 25.00 1.32 24.68 1.32 24.68 0.90 23.60 0.90
                 23.60 1.32 23.28 1.32 23.28 0.90 22.20 0.90 22.20 1.32
                 21.88 1.32 21.88 0.90 20.80 0.90 20.80 1.32 20.48 1.32
                 20.48 0.90 19.40 0.90 19.40 1.32 19.08 1.32 19.08 0.90
                 18.00 0.90 18.00 1.32 17.68 1.32 17.68 0.90 16.60 0.90
                 16.60 1.32 16.28 1.32 16.28 0.90 15.20 0.90 15.20 1.32
                 14.88 1.32 14.88 0.90 13.80 0.90 13.80 1.32 13.48 1.32
                 13.48 0.90 12.40 0.90 12.40 1.32 12.08 1.32 12.08 0.90
                 11.00 0.90 11.00 1.32 10.68 1.32 10.68 0.90 9.60 0.90
                 9.60 1.32 9.28 1.32 9.28 0.90 8.20 0.90 8.20 1.32 7.88 1.32
                 7.88 0.90 6.80 0.90 6.80 1.32 6.48 1.32 6.48 0.90 5.40 0.90
                 5.40 1.32 5.08 1.32 5.08 0.90 4.00 0.90 4.00 1.32 3.68 1.32
                 3.68 0.90 2.60 0.90 2.60 1.32 2.28 1.32 2.28 0.90 1.20 0.90
                 1.20 1.32 0.88 1.32 0.88 0.90 0.00 0.90 0.00 -0.90 34.56 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  34.56 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.34 1.20 4.34
                 1.20 4.86 2.28 4.86 2.28 4.34 2.60 4.34 2.60 4.86 3.68 4.86
                 3.68 4.34 4.00 4.34 4.00 4.86 5.08 4.86 5.08 4.34 5.40 4.34
                 5.40 4.86 6.48 4.86 6.48 4.34 6.80 4.34 6.80 4.86 7.88 4.86
                 7.88 4.34 8.20 4.34 8.20 4.86 9.28 4.86 9.28 4.34 9.60 4.34
                 9.60 4.86 10.68 4.86 10.68 4.34 11.00 4.34 11.00 4.86
                 12.08 4.86 12.08 4.34 12.40 4.34 12.40 4.86 13.48 4.86
                 13.48 4.34 13.80 4.34 13.80 4.86 14.88 4.86 14.88 4.34
                 15.20 4.34 15.20 4.86 16.28 4.86 16.28 4.34 16.60 4.34
                 16.60 4.86 17.68 4.86 17.68 4.34 18.00 4.34 18.00 4.86
                 19.08 4.86 19.08 4.34 19.40 4.34 19.40 4.86 20.48 4.86
                 20.48 4.34 20.80 4.34 20.80 4.86 21.88 4.86 21.88 4.34
                 22.20 4.34 22.20 4.86 23.28 4.86 23.28 4.34 23.60 4.34
                 23.60 4.86 24.68 4.86 24.68 4.34 25.00 4.34 25.00 4.86
                 26.08 4.86 26.08 4.34 26.40 4.34 26.40 4.86 27.48 4.86
                 27.48 4.34 27.80 4.34 27.80 4.86 28.88 4.86 28.88 4.34
                 29.20 4.34 29.20 4.86 30.28 4.86 30.28 4.34 30.60 4.34
                 30.60 4.86 31.68 4.86 31.68 4.34 32.00 4.34 32.00 4.86
                 33.08 4.86 33.08 4.34 33.40 4.34 33.40 4.86 34.56 4.86 ;
        END
    END vdd!
END clkinv_48

MACRO clkinv_4
    CLASS CORE ;
    FOREIGN clkinv_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.84 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.34 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.84  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.30 1.96 1.90 1.96 1.90 3.78 2.98 3.78 2.98 3.28 3.30 3.28
                 3.30 4.10 0.18 4.10 0.18 3.34 0.50 3.34 0.50 3.78 1.58 3.78
                 1.58 3.04 1.44 3.04 1.44 2.72 1.58 2.72 1.58 1.96 0.18 1.96
                 0.18 1.64 3.30 1.64 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  3.84 0.90 2.60 0.90 2.60 1.14 2.28 1.14 2.28 0.90 1.20 0.90
                 1.20 1.14 0.88 1.14 0.88 0.90 0.00 0.90 0.00 -0.90 3.84 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  3.84 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.42 1.20 4.42
                 1.20 4.86 2.28 4.86 2.28 4.42 2.60 4.42 2.60 4.86 3.84 4.86 ;
        END
    END vdd!
END clkinv_4

MACRO clkinv_32
    CLASS CORE ;
    FOREIGN clkinv_32 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 19.93  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.34 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 30.03  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  22.90 1.96 21.50 1.96 21.50 2.72 21.60 2.72 21.60 3.04
                 21.50 3.04 21.50 3.78 22.90 3.78 22.90 4.10 21.18 4.10
                 21.18 1.96 18.70 1.96 18.70 3.78 21.18 3.78 21.18 4.10
                 18.38 4.10 18.38 1.96 15.90 1.96 15.90 3.78 18.38 3.78
                 18.38 4.10 15.58 4.10 15.58 1.96 13.10 1.96 13.10 2.72
                 13.32 2.72 13.32 3.04 13.10 3.04 13.10 3.78 15.58 3.78
                 15.58 4.10 12.78 4.10 12.78 1.96 10.30 1.96 10.30 3.78
                 12.78 3.78 12.78 4.10 9.98 4.10 9.98 1.96 7.50 1.96 7.50 3.78
                 9.98 3.78 9.98 4.10 7.18 4.10 7.18 1.96 4.70 1.96 4.70 3.78
                 7.18 3.78 7.18 4.10 4.38 4.10 4.38 1.96 1.90 1.96 1.90 3.78
                 4.38 3.78 4.38 4.10 0.18 4.10 0.18 3.78 1.58 3.78 1.58 1.96
                 0.18 1.96 0.18 1.64 22.90 1.64 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  23.68 0.90 22.20 0.90 22.20 1.32 21.88 1.32 21.88 0.90
                 20.80 0.90 20.80 1.32 20.48 1.32 20.48 0.90 19.40 0.90
                 19.40 1.32 19.08 1.32 19.08 0.90 18.00 0.90 18.00 1.32
                 17.68 1.32 17.68 0.90 16.60 0.90 16.60 1.32 16.28 1.32
                 16.28 0.90 15.20 0.90 15.20 1.32 14.88 1.32 14.88 0.90
                 13.80 0.90 13.80 1.32 13.48 1.32 13.48 0.90 12.40 0.90
                 12.40 1.32 12.08 1.32 12.08 0.90 11.00 0.90 11.00 1.32
                 10.68 1.32 10.68 0.90 9.60 0.90 9.60 1.32 9.28 1.32 9.28 0.90
                 8.20 0.90 8.20 1.32 7.88 1.32 7.88 0.90 6.80 0.90 6.80 1.32
                 6.48 1.32 6.48 0.90 5.40 0.90 5.40 1.32 5.08 1.32 5.08 0.90
                 4.00 0.90 4.00 1.32 3.68 1.32 3.68 0.90 2.60 0.90 2.60 1.32
                 2.28 1.32 2.28 0.90 1.20 0.90 1.20 1.32 0.88 1.32 0.88 0.90
                 0.00 0.90 0.00 -0.90 23.68 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  23.68 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.42 1.20 4.42
                 1.20 4.86 2.28 4.86 2.28 4.42 2.60 4.42 2.60 4.86 3.68 4.86
                 3.68 4.42 4.00 4.42 4.00 4.86 5.08 4.86 5.08 4.42 5.40 4.42
                 5.40 4.86 6.48 4.86 6.48 4.42 6.80 4.42 6.80 4.86 7.88 4.86
                 7.88 4.42 8.20 4.42 8.20 4.86 9.28 4.86 9.28 4.42 9.60 4.42
                 9.60 4.86 10.68 4.86 10.68 4.42 11.00 4.42 11.00 4.86
                 12.08 4.86 12.08 4.42 12.40 4.42 12.40 4.86 13.48 4.86
                 13.48 4.42 13.80 4.42 13.80 4.86 14.88 4.86 14.88 4.42
                 15.20 4.42 15.20 4.86 16.28 4.86 16.28 4.42 16.60 4.42
                 16.60 4.86 17.68 4.86 17.68 4.42 18.00 4.42 18.00 4.86
                 19.08 4.86 19.08 4.42 19.40 4.42 19.40 4.86 20.48 4.86
                 20.48 4.42 20.80 4.42 20.80 4.86 21.88 4.86 21.88 4.42
                 22.20 4.42 22.20 4.86 23.68 4.86 ;
        END
    END vdd!
END clkinv_32

MACRO clkinv_3
    CLASS CORE ;
    FOREIGN clkinv_3 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.20 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.87  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.34 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.32  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.90 4.38 1.58 4.38 1.58 3.88 0.50 3.88 0.50 4.38 0.18 4.38
                 0.18 3.34 0.50 3.34 0.50 3.56 1.58 3.56 1.58 3.04 1.44 3.04
                 1.44 2.72 1.58 2.72 1.58 1.96 0.18 1.96 0.18 1.64 1.90 1.64 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  3.20 0.90 2.60 0.90 2.60 2.18 2.28 2.18 2.28 0.90 1.20 0.90
                 1.20 1.14 0.88 1.14 0.88 0.90 0.00 0.90 0.00 -0.90 3.20 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  3.20 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.34 1.20 4.34
                 1.20 4.86 2.28 4.86 2.28 3.28 2.60 3.28 2.60 4.86 3.20 4.86 ;
        END
    END vdd!
END clkinv_3

MACRO clkinv_24
    CLASS CORE ;
    FOREIGN clkinv_24 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 17.92 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 14.95  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.34 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 22.84  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  17.30 1.96 15.90 1.96 15.90 3.56 16.98 3.56 16.98 3.34
                 17.30 3.34 17.30 4.38 16.98 4.38 16.98 3.88 15.90 3.88
                 15.90 4.38 15.58 4.38 15.58 3.22 15.52 3.22 15.52 2.72
                 15.58 2.72 15.58 1.96 14.50 1.96 14.50 3.56 15.58 3.56
                 15.58 3.88 14.50 3.88 14.50 4.38 14.18 4.38 14.18 1.96
                 11.70 1.96 11.70 3.56 12.78 3.56 12.78 3.34 13.10 3.34
                 13.10 3.56 14.18 3.56 14.18 3.88 13.10 3.88 13.10 4.38
                 12.78 4.38 12.78 3.88 11.70 3.88 11.70 4.38 11.38 4.38
                 11.38 1.96 10.30 1.96 10.30 3.56 11.38 3.56 11.38 3.88
                 10.30 3.88 10.30 4.38 9.98 4.38 9.98 1.96 7.50 1.96 7.50 3.56
                 8.58 3.56 8.58 3.34 8.90 3.34 8.90 3.56 9.98 3.56 9.98 3.88
                 8.90 3.88 8.90 4.38 8.58 4.38 8.58 3.88 7.50 3.88 7.50 4.38
                 7.18 4.38 7.18 1.96 6.10 1.96 6.10 3.56 7.18 3.56 7.18 3.88
                 6.10 3.88 6.10 4.38 5.78 4.38 5.78 1.96 3.30 1.96 3.30 3.56
                 4.38 3.56 4.38 3.34 4.70 3.34 4.70 3.56 5.78 3.56 5.78 3.88
                 4.70 3.88 4.70 4.38 4.38 4.38 4.38 3.88 3.30 3.88 3.30 4.38
                 2.98 4.38 2.98 1.96 1.90 1.96 1.90 3.56 2.98 3.56 2.98 3.88
                 1.90 3.88 1.90 4.38 1.58 4.38 1.58 3.88 0.50 3.88 0.50 4.38
                 0.18 4.38 0.18 3.34 0.50 3.34 0.50 3.56 1.58 3.56 1.58 1.96
                 0.18 1.96 0.18 1.64 17.30 1.64 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  17.92 0.90 16.60 0.90 16.60 1.32 16.28 1.32 16.28 0.90
                 15.20 0.90 15.20 1.32 14.88 1.32 14.88 0.90 13.80 0.90
                 13.80 1.32 13.48 1.32 13.48 0.90 12.40 0.90 12.40 1.32
                 12.08 1.32 12.08 0.90 11.00 0.90 11.00 1.32 10.68 1.32
                 10.68 0.90 9.60 0.90 9.60 1.32 9.28 1.32 9.28 0.90 8.20 0.90
                 8.20 1.32 7.88 1.32 7.88 0.90 6.80 0.90 6.80 1.32 6.48 1.32
                 6.48 0.90 5.40 0.90 5.40 1.32 5.08 1.32 5.08 0.90 4.00 0.90
                 4.00 1.32 3.68 1.32 3.68 0.90 2.60 0.90 2.60 1.32 2.28 1.32
                 2.28 0.90 1.20 0.90 1.20 1.32 0.88 1.32 0.88 0.90 0.00 0.90
                 0.00 -0.90 17.92 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  17.92 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.34 1.20 4.34
                 1.20 4.86 2.28 4.86 2.28 4.34 2.60 4.34 2.60 4.86 3.68 4.86
                 3.68 4.34 4.00 4.34 4.00 4.86 5.08 4.86 5.08 4.34 5.40 4.34
                 5.40 4.86 6.48 4.86 6.48 4.34 6.80 4.34 6.80 4.86 7.88 4.86
                 7.88 4.34 8.20 4.34 8.20 4.86 9.28 4.86 9.28 4.34 9.60 4.34
                 9.60 4.86 10.68 4.86 10.68 4.34 11.00 4.34 11.00 4.86
                 12.08 4.86 12.08 4.34 12.40 4.34 12.40 4.86 13.48 4.86
                 13.48 4.34 13.80 4.34 13.80 4.86 14.88 4.86 14.88 4.34
                 15.20 4.34 15.20 4.86 16.28 4.86 16.28 4.34 16.60 4.34
                 16.60 4.86 17.92 4.86 ;
        END
    END vdd!
END clkinv_24

MACRO clkinv_20
    CLASS CORE ;
    FOREIGN clkinv_20 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.72 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 12.46  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.34 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 19.24  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  14.50 1.96 13.10 1.96 13.10 2.72 13.28 2.72 13.28 3.04
                 13.10 3.04 13.10 3.58 14.50 3.58 14.50 4.54 14.18 4.54
                 14.18 3.90 13.10 3.90 13.10 4.54 12.78 4.54 12.78 1.96
                 8.90 1.96 8.90 3.58 12.78 3.58 12.78 3.90 11.70 3.90
                 11.70 4.54 11.38 4.54 11.38 3.90 10.30 3.90 10.30 4.54
                 9.98 4.54 9.98 3.90 8.90 3.90 8.90 4.54 8.58 4.54 8.58 1.96
                 6.10 1.96 6.10 3.58 8.58 3.58 8.58 3.90 7.50 3.90 7.50 4.54
                 7.18 4.54 7.18 3.90 6.10 3.90 6.10 4.54 5.78 4.54 5.78 1.96
                 1.90 1.96 1.90 3.58 5.78 3.58 5.78 3.90 4.70 3.90 4.70 4.54
                 4.38 4.54 4.38 3.90 3.30 3.90 3.30 4.54 2.98 4.54 2.98 3.90
                 1.90 3.90 1.90 4.54 1.58 4.54 1.58 3.90 0.50 3.90 0.50 4.54
                 0.18 4.54 0.18 3.58 1.58 3.58 1.58 1.96 0.18 1.96 0.18 1.64
                 14.50 1.64 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  14.72 0.90 13.80 0.90 13.80 1.32 13.48 1.32 13.48 0.90
                 12.40 0.90 12.40 1.32 12.08 1.32 12.08 0.90 11.00 0.90
                 11.00 1.32 10.68 1.32 10.68 0.90 9.60 0.90 9.60 1.32 9.28 1.32
                 9.28 0.90 8.20 0.90 8.20 1.32 7.88 1.32 7.88 0.90 6.80 0.90
                 6.80 1.32 6.48 1.32 6.48 0.90 5.40 0.90 5.40 1.32 5.08 1.32
                 5.08 0.90 4.00 0.90 4.00 1.32 3.68 1.32 3.68 0.90 2.60 0.90
                 2.60 1.32 2.28 1.32 2.28 0.90 1.20 0.90 1.20 1.32 0.88 1.32
                 0.88 0.90 0.00 0.90 0.00 -0.90 14.72 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  14.72 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 2.28 4.86 2.28 4.22 2.60 4.22 2.60 4.86 3.68 4.86
                 3.68 4.22 4.00 4.22 4.00 4.86 5.08 4.86 5.08 4.22 5.40 4.22
                 5.40 4.86 6.48 4.86 6.48 4.22 6.80 4.22 6.80 4.86 7.88 4.86
                 7.88 4.22 8.20 4.22 8.20 4.86 9.28 4.86 9.28 4.22 9.60 4.22
                 9.60 4.86 10.68 4.86 10.68 4.22 11.00 4.22 11.00 4.86
                 12.08 4.86 12.08 4.22 12.40 4.22 12.40 4.86 13.48 4.86
                 13.48 4.22 13.80 4.22 13.80 4.86 14.72 4.86 ;
        END
    END vdd!
END clkinv_20

MACRO clkinv_2
    CLASS CORE ;
    FOREIGN clkinv_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.56 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.25  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.34 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.04  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.90 4.32 1.58 4.32 1.58 4.04 0.50 4.04 0.50 4.32 0.18 4.32
                 0.18 3.44 0.50 3.44 0.50 3.72 1.58 3.72 1.58 3.04 1.44 3.04
                 1.44 2.72 1.58 2.72 1.58 1.96 0.18 1.96 0.18 1.64 1.90 1.64 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  2.56 0.90 1.20 0.90 1.20 1.15 0.88 1.15 0.88 0.90 0.00 0.90
                 0.00 -0.90 2.56 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  2.56 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.42 1.20 4.42
                 1.20 4.86 2.56 4.86 ;
        END
    END vdd!
END clkinv_2

MACRO clkinv_16
    CLASS CORE ;
    FOREIGN clkinv_16 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.16 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 9.96  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.34 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 15.64  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  11.70 1.96 10.30 1.96 10.30 3.78 11.70 3.78 11.70 4.10
                 9.98 4.10 9.98 3.04 9.76 3.04 9.76 2.72 9.98 2.72 9.98 1.96
                 7.50 1.96 7.50 3.78 9.98 3.78 9.98 4.10 7.18 4.10 7.18 1.96
                 4.70 1.96 4.70 3.78 7.18 3.78 7.18 4.10 4.38 4.10 4.38 1.96
                 1.90 1.96 1.90 3.78 4.38 3.78 4.38 4.10 0.18 4.10 0.18 3.78
                 1.58 3.78 1.58 1.96 0.18 1.96 0.18 1.64 11.70 1.64 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  12.16 0.90 11.00 0.90 11.00 1.32 10.68 1.32 10.68 0.90
                 9.60 0.90 9.60 1.32 9.28 1.32 9.28 0.90 8.20 0.90 8.20 1.32
                 7.88 1.32 7.88 0.90 6.80 0.90 6.80 1.32 6.48 1.32 6.48 0.90
                 5.40 0.90 5.40 1.32 5.08 1.32 5.08 0.90 4.00 0.90 4.00 1.32
                 3.68 1.32 3.68 0.90 2.60 0.90 2.60 1.32 2.28 1.32 2.28 0.90
                 1.20 0.90 1.20 1.32 0.88 1.32 0.88 0.90 0.00 0.90 0.00 -0.90
                 12.16 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  12.16 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.42 1.20 4.42
                 1.20 4.86 2.28 4.86 2.28 4.42 2.60 4.42 2.60 4.86 3.68 4.86
                 3.68 4.42 4.00 4.42 4.00 4.86 5.08 4.86 5.08 4.42 5.40 4.42
                 5.40 4.86 6.48 4.86 6.48 4.42 6.80 4.42 6.80 4.86 7.88 4.86
                 7.88 4.42 8.20 4.42 8.20 4.86 9.28 4.86 9.28 4.42 9.60 4.42
                 9.60 4.86 10.68 4.86 10.68 4.42 11.00 4.42 11.00 4.86
                 12.16 4.86 ;
        END
    END vdd!
END clkinv_16

MACRO clkinv_12
    CLASS CORE ;
    FOREIGN clkinv_12 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.60 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 7.47  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.34 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 12.04  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.90 1.96 7.50 1.96 7.50 2.72 7.52 2.72 7.52 3.04 7.50 3.04
                 7.50 3.56 8.58 3.56 8.58 3.34 8.90 3.34 8.90 4.38 8.58 4.38
                 8.58 3.88 7.50 3.88 7.50 4.38 7.18 4.38 7.18 1.96 6.10 1.96
                 6.10 3.56 7.18 3.56 7.18 3.88 6.10 3.88 6.10 4.38 5.78 4.38
                 5.78 1.96 3.30 1.96 3.30 3.56 4.38 3.56 4.38 3.34 4.70 3.34
                 4.70 3.56 5.78 3.56 5.78 3.88 4.70 3.88 4.70 4.38 4.38 4.38
                 4.38 3.88 3.30 3.88 3.30 4.38 2.98 4.38 2.98 1.96 1.90 1.96
                 1.90 3.56 2.98 3.56 2.98 3.88 1.90 3.88 1.90 4.38 1.58 4.38
                 1.58 3.88 0.50 3.88 0.50 4.38 0.18 4.38 0.18 3.34 0.50 3.34
                 0.50 3.56 1.58 3.56 1.58 1.96 0.18 1.96 0.18 1.64 8.90 1.64 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  9.60 0.90 8.20 0.90 8.20 1.32 7.88 1.32 7.88 0.90 6.80 0.90
                 6.80 1.32 6.48 1.32 6.48 0.90 5.40 0.90 5.40 1.32 5.08 1.32
                 5.08 0.90 4.00 0.90 4.00 1.32 3.68 1.32 3.68 0.90 2.60 0.90
                 2.60 1.32 2.28 1.32 2.28 0.90 1.20 0.90 1.20 1.32 0.88 1.32
                 0.88 0.90 0.00 0.90 0.00 -0.90 9.60 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  9.60 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.34 1.20 4.34
                 1.20 4.86 2.28 4.86 2.28 4.34 2.60 4.34 2.60 4.86 3.68 4.86
                 3.68 4.34 4.00 4.34 4.00 4.86 5.08 4.86 5.08 4.34 5.40 4.34
                 5.40 4.86 6.48 4.86 6.48 4.34 6.80 4.34 6.80 4.86 7.88 4.86
                 7.88 4.34 8.20 4.34 8.20 4.86 9.60 4.86 ;
        END
    END vdd!
END clkinv_12

MACRO clkinv_10
    CLASS CORE ;
    FOREIGN clkinv_10 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 6.23  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.34 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 10.24  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.50 1.96 6.10 1.96 6.10 2.72 6.24 2.72 6.24 3.04 6.10 3.04
                 6.10 3.58 7.50 3.58 7.50 4.54 7.18 4.54 7.18 3.90 6.10 3.90
                 6.10 4.54 5.78 4.54 5.78 1.96 1.90 1.96 1.90 3.58 5.78 3.58
                 5.78 3.90 4.70 3.90 4.70 4.54 4.38 4.54 4.38 3.90 3.30 3.90
                 3.30 4.54 2.98 4.54 2.98 3.90 1.90 3.90 1.90 4.54 1.58 4.54
                 1.58 3.90 0.50 3.90 0.50 4.54 0.18 4.54 0.18 3.58 1.58 3.58
                 1.58 1.96 0.18 1.96 0.18 1.64 7.50 1.64 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 0.90 6.80 0.90 6.80 1.32 6.48 1.32 6.48 0.90 5.40 0.90
                 5.40 1.32 5.08 1.32 5.08 0.90 4.00 0.90 4.00 1.32 3.68 1.32
                 3.68 0.90 2.60 0.90 2.60 1.32 2.28 1.32 2.28 0.90 1.20 0.90
                 1.20 1.32 0.88 1.32 0.88 0.90 0.00 0.90 0.00 -0.90 7.68 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 2.28 4.86 2.28 4.22 2.60 4.22 2.60 4.86 3.68 4.86
                 3.68 4.22 4.00 4.22 4.00 4.86 5.08 4.86 5.08 4.22 5.40 4.22
                 5.40 4.86 6.48 4.86 6.48 4.22 6.80 4.22 6.80 4.86 7.68 4.86 ;
        END
    END vdd!
END clkinv_10

MACRO clkinv_1
    CLASS CORE ;
    FOREIGN clkinv_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 1.92 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.62  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.48 2.62 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.51  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.76 3.78 1.44 3.78 1.44 4.54 1.12 4.54 1.12 3.46 1.44 3.46
                 1.44 2.04 1.12 2.04 1.12 1.72 1.76 1.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  1.92 0.90 0.74 0.90 0.74 1.40 0.42 1.40 0.42 0.90 0.00 0.90
                 0.00 -0.90 1.92 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  1.92 6.66 0.00 6.66 0.00 4.86 0.42 4.86 0.42 3.56 0.74 3.56
                 0.74 4.86 1.92 4.86 ;
        END
    END vdd!
END clkinv_1

MACRO clkinv_0
    CLASS CORE ;
    FOREIGN clkinv_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 1.92 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.54  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.48 2.62 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.31  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  1.76 3.78 1.44 3.78 1.44 4.34 1.12 4.34 1.12 3.46 1.44 3.46
                 1.44 2.11 1.12 2.11 1.12 1.79 1.76 1.79 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  1.92 0.90 0.74 0.90 0.74 1.62 0.42 1.62 0.42 0.90 0.00 0.90
                 0.00 -0.90 1.92 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  1.92 6.66 0.00 6.66 0.00 4.86 0.42 4.86 0.42 3.56 0.74 3.56
                 0.74 4.86 1.92 4.86 ;
        END
    END vdd!
END clkinv_0

MACRO clkbuf_8
    CLASS CORE ;
    FOREIGN clkbuf_8 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.80 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 4.22  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.58 2.43 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 8.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.38 1.55 12.00 1.55 12.00 3.76 12.38 3.76 12.38 4.08
                 11.68 4.08 11.68 1.55 8.46 1.55 8.46 3.76 11.68 3.76
                 11.68 4.08 6.46 4.08 6.46 3.76 8.14 3.76 8.14 1.55 6.46 1.55
                 6.46 1.23 12.38 1.23 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 12.80 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 12.80 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  7.77 3.09 6.10 3.09 6.10 4.16 5.78 4.16 5.78 1.61 1.90 1.61
                 1.90 3.84 5.78 3.84 5.78 4.16 0.18 4.16 0.18 3.84 1.58 3.84
                 1.58 1.61 0.18 1.61 0.18 1.29 6.10 1.29 6.10 2.77 7.77 2.77 ;
    END
END clkbuf_8

MACRO clkbuf_64
    CLASS CORE ;
    FOREIGN clkbuf_64 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 91.52 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 33.75  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.58 2.43 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 57.12  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  90.78 4.08 90.46 4.08 90.46 3.04 90.40 3.04 90.40 2.72
                 90.46 2.72 90.46 1.54 85.19 1.54 85.19 3.76 90.46 3.76
                 90.46 4.08 84.87 4.08 84.87 1.54 79.58 1.54 79.58 3.76
                 84.87 3.76 84.87 4.08 79.26 4.08 79.26 1.54 73.98 1.54
                 73.98 3.76 79.26 3.76 79.26 4.08 73.66 4.08 73.66 1.54
                 68.38 1.54 68.38 3.76 73.66 3.76 73.66 4.08 68.06 4.08
                 68.06 1.54 62.78 1.54 62.78 3.76 68.06 3.76 68.06 4.08
                 62.46 4.08 62.46 1.54 57.18 1.54 57.18 3.76 62.46 3.76
                 62.46 4.08 56.86 4.08 56.86 1.54 51.58 1.54 51.58 3.76
                 56.86 3.76 56.86 4.08 51.26 4.08 51.26 1.54 47.67 1.54
                 47.67 3.76 51.26 3.76 51.26 4.08 45.66 4.08 45.66 3.76
                 47.35 3.76 47.35 1.54 45.66 1.54 45.66 1.22 90.78 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 91.52 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 91.52 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  46.97 3.08 45.30 3.08 45.30 4.16 44.98 4.16 44.98 1.61
                 39.70 1.61 39.70 3.84 44.98 3.84 44.98 4.16 39.38 4.16
                 39.38 1.61 34.10 1.61 34.10 3.84 39.38 3.84 39.38 4.16
                 33.78 4.16 33.78 1.61 28.50 1.61 28.50 3.84 33.78 3.84
                 33.78 4.16 28.18 4.16 28.18 1.61 22.90 1.61 22.90 3.84
                 28.18 3.84 28.18 4.16 22.58 4.16 22.58 1.61 17.30 1.61
                 17.30 3.84 22.58 3.84 22.58 4.16 16.98 4.16 16.98 1.61
                 11.70 1.61 11.70 3.84 16.98 3.84 16.98 4.16 11.38 4.16
                 11.38 1.61 6.10 1.61 6.10 3.84 11.38 3.84 11.38 4.16 5.78 4.16
                 5.78 1.61 1.90 1.61 1.90 3.84 5.78 3.84 5.78 4.16 0.18 4.16
                 0.18 3.84 1.58 3.84 1.58 1.61 0.18 1.61 0.18 1.29 45.30 1.29
                 45.30 2.76 46.97 2.76 ;
    END
END clkbuf_64

MACRO clkbuf_6
    CLASS CORE ;
    FOREIGN clkbuf_6 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.24 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.16  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.58 2.43 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.45  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.58 1.55 9.44 1.55 9.44 3.76 9.58 3.76 9.58 4.08 5.06 4.08
                 5.06 3.76 9.12 3.76 9.12 1.55 5.06 1.55 5.06 1.23 9.58 1.23 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 10.24 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 10.24 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  6.37 3.09 4.70 3.09 4.70 4.16 4.38 4.16 4.38 1.61 1.90 1.61
                 1.90 3.84 4.38 3.84 4.38 4.16 0.18 4.16 0.18 3.84 1.58 3.84
                 1.58 1.61 0.18 1.61 0.18 1.29 4.70 1.29 4.70 2.77 6.37 2.77 ;
    END
END clkbuf_6

MACRO clkbuf_48
    CLASS CORE ;
    FOREIGN clkbuf_48 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 69.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 25.32  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.58 2.43 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 43.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  68.38 4.54 68.06 4.54 68.06 3.04 68.00 3.04 68.00 2.72
                 68.06 2.72 68.06 1.55 62.78 1.55 62.78 4.22 68.06 4.22
                 68.06 4.54 62.46 4.54 62.46 1.55 57.18 1.55 57.18 4.22
                 62.46 4.22 62.46 4.54 56.86 4.54 56.86 1.55 51.58 1.55
                 51.58 4.22 56.86 4.22 56.86 4.54 51.26 4.54 51.26 1.55
                 45.98 1.55 45.98 4.22 51.26 4.22 51.26 4.54 45.66 4.54
                 45.66 1.55 40.38 1.55 40.38 4.22 45.66 4.22 45.66 4.54
                 40.06 4.54 40.06 1.55 36.47 1.55 36.47 4.22 40.06 4.22
                 40.06 4.54 34.46 4.54 34.46 4.22 36.15 4.22 36.15 1.55
                 34.46 1.55 34.46 1.23 68.38 1.23 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 69.12 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 69.12 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  35.77 3.08 34.10 3.08 34.10 4.16 33.78 4.16 33.78 1.61
                 28.50 1.61 28.50 3.84 33.78 3.84 33.78 4.16 28.18 4.16
                 28.18 1.61 22.90 1.61 22.90 3.84 28.18 3.84 28.18 4.16
                 22.58 4.16 22.58 1.61 17.30 1.61 17.30 3.84 22.58 3.84
                 22.58 4.16 16.98 4.16 16.98 1.61 11.70 1.61 11.70 3.84
                 16.98 3.84 16.98 4.16 11.38 4.16 11.38 1.61 6.10 1.61
                 6.10 3.84 11.38 3.84 11.38 4.16 5.78 4.16 5.78 1.61 1.76 1.61
                 1.76 3.84 5.78 3.84 5.78 4.16 0.18 4.16 0.18 3.84 1.44 3.84
                 1.44 1.61 0.18 1.61 0.18 1.29 34.10 1.29 34.10 2.75 35.77 2.75 ;
    END
END clkbuf_48

MACRO clkbuf_4
    CLASS CORE ;
    FOREIGN clkbuf_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.04 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.11  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.58 2.43 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.70  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  6.88 4.08 3.66 4.08 3.66 3.76 6.56 3.76 6.56 1.55 3.66 1.55
                 3.66 1.23 6.88 1.23 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 7.04 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 7.04 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.97 3.09 3.30 3.09 3.30 4.16 0.18 4.16 0.18 3.84 2.98 3.84
                 2.98 1.61 0.18 1.61 0.18 1.29 3.30 1.29 3.30 2.77 4.97 2.77 ;
    END
END clkbuf_4

MACRO clkbuf_32
    CLASS CORE ;
    FOREIGN clkbuf_32 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 46.72 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 16.93  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.58 2.43 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 29.16  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  45.98 4.08 45.66 4.08 45.66 3.04 45.60 3.04 45.60 2.72
                 45.66 2.72 45.66 1.54 40.38 1.54 40.38 3.76 45.66 3.76
                 45.66 4.08 40.06 4.08 40.06 1.54 34.78 1.54 34.78 3.76
                 40.06 3.76 40.06 4.08 34.46 4.08 34.46 1.54 29.18 1.54
                 29.18 3.76 34.46 3.76 34.46 4.08 28.86 4.08 28.86 1.54
                 25.27 1.54 25.27 3.76 28.86 3.76 28.86 4.08 23.26 4.08
                 23.26 3.76 24.95 3.76 24.95 1.54 23.26 1.54 23.26 1.22
                 45.98 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 46.72 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 46.72 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  24.57 3.09 22.90 3.09 22.90 4.15 22.58 4.15 22.58 1.61
                 17.30 1.61 17.30 3.83 22.58 3.83 22.58 4.15 16.98 4.15
                 16.98 1.61 11.70 1.61 11.70 3.83 16.98 3.83 16.98 4.15
                 11.38 4.15 11.38 1.61 6.10 1.61 6.10 3.83 11.38 3.83
                 11.38 4.15 5.78 4.15 5.78 1.61 1.76 1.61 1.76 3.83 5.78 3.83
                 5.78 4.15 0.18 4.15 0.18 3.83 1.44 3.83 1.44 1.61 0.18 1.61
                 0.18 1.29 22.90 1.29 22.90 2.77 24.57 2.77 ;
    END
END clkbuf_32

MACRO clkbuf_3
    CLASS CORE ;
    FOREIGN clkbuf_3 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.48 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.05  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.58 2.43 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.96  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.32 4.08 2.26 4.08 2.26 3.76 4.00 3.76 4.00 1.55 2.26 1.55
                 2.26 1.23 4.32 1.23 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 4.48 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 4.48 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  3.57 3.09 1.90 3.09 1.90 4.16 0.18 4.16 0.18 3.84 1.58 3.84
                 1.58 1.61 0.18 1.61 0.18 1.29 1.90 1.29 1.90 2.77 3.57 2.77 ;
    END
END clkbuf_3

MACRO clkbuf_24
    CLASS CORE ;
    FOREIGN clkbuf_24 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 35.20 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 12.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.58 2.43 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 22.18  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  34.78 1.55 34.40 1.55 34.40 3.76 34.78 3.76 34.78 4.08
                 34.08 4.08 34.08 1.55 29.18 1.55 29.18 3.76 34.08 3.76
                 34.08 4.08 28.86 4.08 28.86 1.55 23.58 1.55 23.58 3.76
                 28.86 3.76 28.86 4.08 23.26 4.08 23.26 1.55 19.67 1.55
                 19.67 3.76 23.26 3.76 23.26 4.08 17.66 4.08 17.66 3.76
                 19.35 3.76 19.35 1.55 17.66 1.55 17.66 1.23 34.78 1.23 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 35.20 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 35.20 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  18.97 3.09 17.30 3.09 17.30 4.16 16.98 4.16 16.98 1.61
                 11.70 1.61 11.70 3.84 16.98 3.84 16.98 4.16 11.38 4.16
                 11.38 1.61 6.10 1.61 6.10 3.84 11.38 3.84 11.38 4.16 0.18 4.16
                 0.18 3.84 5.78 3.84 5.78 1.61 0.18 1.61 0.18 1.29 17.30 1.29
                 17.30 2.77 18.97 2.77 ;
    END
END clkbuf_24

MACRO clkbuf_20
    CLASS CORE ;
    FOREIGN clkbuf_20 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 29.44 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 10.55  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.58 2.43 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 18.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  29.18 1.55 28.00 1.55 28.00 3.76 29.18 3.76 29.18 4.08
                 27.68 4.08 27.68 1.55 22.18 1.55 22.18 3.76 27.68 3.76
                 27.68 4.08 21.86 4.08 21.86 1.55 16.87 1.55 16.87 3.76
                 21.86 3.76 21.86 4.08 14.86 4.08 14.86 3.76 16.55 3.76
                 16.55 1.55 14.86 1.55 14.86 1.23 29.18 1.23 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 29.44 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 29.44 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  16.17 3.09 14.50 3.09 14.50 4.16 14.18 4.16 14.18 1.61
                 8.90 1.61 8.90 3.84 14.18 3.84 14.18 4.16 8.58 4.16 8.58 1.61
                 3.30 1.61 3.30 3.84 8.58 3.84 8.58 4.16 0.18 4.16 0.18 3.84
                 2.98 3.84 2.98 1.61 0.18 1.61 0.18 1.29 14.50 1.29 14.50 2.77
                 16.17 2.77 ;
    END
END clkbuf_20

MACRO clkbuf_2
    CLASS CORE ;
    FOREIGN clkbuf_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.58  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.58 2.43 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.23  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.96 4.08 3.21 4.08 3.21 3.76 4.64 3.76 4.64 1.55 3.22 1.55
                 3.22 1.23 4.96 1.23 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 5.12 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 5.12 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  3.81 3.09 1.90 3.09 1.90 4.16 0.18 4.16 0.18 3.84 1.58 3.84
                 1.58 1.61 0.18 1.61 0.18 1.29 1.90 1.29 1.90 2.77 3.81 2.77 ;
    END
END clkbuf_2

MACRO clkbuf_16
    CLASS CORE ;
    FOREIGN clkbuf_16 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 24.32 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 8.44  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.58 2.43 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 15.19  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  23.59 1.55 21.60 1.55 21.60 3.76 23.59 3.76 23.59 4.08
                 21.28 4.08 21.28 1.55 14.08 1.55 14.08 3.76 21.28 3.76
                 21.28 4.08 12.07 4.08 12.07 3.76 13.76 3.76 13.76 1.55
                 12.07 1.55 12.07 1.23 23.59 1.23 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 24.32 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 24.32 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  13.38 3.09 11.71 3.09 11.71 4.16 11.39 4.16 11.39 1.61
                 6.11 1.61 6.11 3.84 11.39 3.84 11.39 4.16 5.79 4.16 5.79 1.61
                 1.87 1.61 1.87 3.84 5.79 3.84 5.79 4.16 0.19 4.16 0.19 3.84
                 1.55 3.84 1.55 1.61 0.19 1.61 0.19 1.29 11.71 1.29 11.71 2.77
                 13.38 2.77 ;
    END
END clkbuf_16

MACRO clkbuf_12
    CLASS CORE ;
    FOREIGN clkbuf_12 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.56 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 6.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.66 2.43 1.20 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 11.69  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  18.06 1.55 17.76 1.55 17.76 3.76 18.06 3.76 18.06 4.08
                 17.44 4.08 17.44 1.55 11.35 1.55 11.35 3.76 17.44 3.76
                 17.44 4.08 9.34 4.08 9.34 3.76 11.03 3.76 11.03 1.55 9.34 1.55
                 9.34 1.23 18.06 1.23 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 18.56 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 18.56 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  10.65 3.09 8.98 3.09 8.98 4.16 8.66 4.16 8.66 1.61 3.38 1.61
                 3.38 3.84 8.66 3.84 8.66 4.16 0.26 4.16 0.26 3.84 3.06 3.84
                 3.06 1.61 0.26 1.61 0.26 1.29 8.98 1.29 8.98 2.77 10.65 2.77 ;
    END
END clkbuf_12

MACRO clkbuf_10
    CLASS CORE ;
    FOREIGN clkbuf_10 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.36 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 5.27  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.58 2.43 1.12 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 9.95  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  15.18 1.55 14.56 1.55 14.56 3.76 15.18 3.76 15.18 4.08
                 14.24 4.08 14.24 1.55 9.86 1.55 9.86 3.76 14.24 3.76
                 14.24 4.08 7.86 4.08 7.86 3.76 9.54 3.76 9.54 1.55 7.86 1.55
                 7.86 1.23 15.18 1.23 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 15.36 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 15.36 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  9.17 3.09 7.50 3.09 7.50 4.16 7.18 4.16 7.18 1.61 1.90 1.61
                 1.90 3.84 7.18 3.84 7.18 4.16 0.18 4.16 0.18 3.84 1.58 3.84
                 1.58 1.61 0.18 1.61 0.18 1.29 7.50 1.29 7.50 2.77 9.17 2.77 ;
    END
END clkbuf_10

MACRO clkbuf_1
    CLASS CORE ;
    FOREIGN clkbuf_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.56 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.53  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.44 2.41 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.48  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  2.40 4.15 1.82 4.15 1.82 3.83 2.08 3.83 2.08 1.57 1.82 1.57
                 1.82 1.25 2.40 1.25 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  2.56 0.90 1.28 0.90 1.28 1.61 0.96 1.61 0.96 0.90 0.00 0.90
                 0.00 -0.90 2.56 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  2.56 6.66 0.00 6.66 0.00 4.86 0.98 4.86 0.98 4.34 1.30 4.34
                 1.30 4.86 2.56 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  1.72 3.09 0.48 3.09 0.48 3.83 0.50 3.83 0.50 4.15 0.16 4.15
                 0.16 1.29 0.50 1.29 0.50 1.61 0.48 1.61 0.48 2.77 1.72 2.77 ;
    END
END clkbuf_1

MACRO clkbuf_0
    CLASS CORE ;
    FOREIGN clkbuf_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.56 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.52  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.00 1.12 2.64 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.28  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  2.40 4.16 1.82 4.16 1.82 3.84 2.08 3.84 2.08 1.58 1.82 1.58
                 1.82 1.26 2.40 1.26 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 2.56 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 2.56 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  1.72 3.41 0.48 3.41 0.48 3.84 0.74 3.84 0.74 4.16 0.16 4.16
                 0.16 1.26 0.74 1.26 0.74 1.58 0.48 1.58 0.48 3.09 1.72 3.09 ;
    END
END clkbuf_0

MACRO busholden1
    CLASS CORE ;
    FOREIGN busholden1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.76 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INOUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.32  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  5.60 3.68 5.36 3.68 5.36 4.54 5.04 4.54 5.04 3.36 5.28 3.36
                 5.28 2.08 4.34 2.08 4.34 2.18 3.27 2.18 3.27 2.43 2.95 2.43
                 2.95 1.86 4.02 1.86 4.02 1.76 5.60 1.76 ;
        END
    END a
    PIN en
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.32  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.24 2.08 1.76 2.69 ;
        END
    END en
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  5.76 0.90 4.66 0.90 4.66 1.32 4.34 1.32 4.34 0.90 0.00 0.90
                 0.00 -0.90 5.76 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.76 6.66 0.00 6.66 0.00 4.86 2.96 4.86 2.96 4.29 3.28 4.29
                 3.28 4.86 4.34 4.86 4.34 3.56 4.66 3.56 4.66 4.86 5.76 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.96 2.91 3.98 2.91 3.98 3.33 0.50 3.33 0.50 4.33 0.18 4.33
                 0.18 3.01 0.58 3.01 0.58 1.22 3.70 1.22 3.70 1.54 0.90 1.54
                 0.90 3.01 3.66 3.01 3.66 2.59 4.96 2.59 ;
        POLYGON  3.98 4.54 3.66 4.54 3.66 3.97 1.20 3.97 1.20 4.54 0.88 4.54
                 0.88 3.65 3.98 3.65 ;
    END
END busholden1

MACRO busholden0
    CLASS CORE ;
    FOREIGN busholden0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.76 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INOUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.13  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  5.60 3.90 3.41 3.90 3.41 3.68 2.08 3.68 2.08 2.94 2.46 2.94
                 2.46 3.36 3.73 3.36 3.73 3.58 5.28 3.58 5.28 1.70 5.04 1.70
                 5.04 1.38 5.60 1.38 ;
        END
    END a
    PIN en
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.13  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.62 1.76 3.26 ;
        END
    END en
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  5.76 0.90 4.66 0.90 4.66 1.32 4.34 1.32 4.34 0.90 0.00 0.90
                 0.00 -0.90 5.76 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.76 6.66 0.00 6.66 0.00 4.86 4.34 4.86 4.34 4.30 4.66 4.30
                 4.66 4.86 5.76 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.96 2.66 3.73 2.66 3.73 2.22 1.12 2.22 1.12 4.22 3.64 4.22
                 3.64 4.54 0.52 4.54 0.52 4.22 0.80 4.22 0.80 2.22 0.18 2.22
                 0.18 1.22 0.50 1.22 0.50 1.90 4.05 1.90 4.05 2.34 4.96 2.34 ;
        RECT  0.88 1.22 3.98 1.54 ;
    END
END busholden0

MACRO bushold
    CLASS CORE ;
    FOREIGN bushold 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.56 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INOUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  2.36 3.90 2.14 3.90 2.14 4.54 1.82 4.54 1.82 3.58 2.04 3.58
                 2.04 2.27 1.12 2.27 1.12 2.45 0.80 2.45 0.80 1.94 2.04 1.94
                 2.04 1.54 1.82 1.54 1.82 1.22 2.36 1.22 ;
        END
    END a
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  2.56 0.90 1.32 0.90 1.32 1.54 1.00 1.54 1.00 0.90 0.00 0.90
                 0.00 -0.90 2.56 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  2.56 6.66 0.00 6.66 0.00 4.86 0.98 4.86 0.98 3.58 1.30 3.58
                 1.30 4.86 2.56 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  1.72 3.09 0.48 3.09 0.48 3.58 0.50 3.58 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 2.77 1.40 2.77
                 1.40 2.62 1.72 2.62 ;
    END
END bushold

MACRO buf_8
    CLASS CORE ;
    FOREIGN buf_8 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.47 0.82 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.29  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.96 4.54 1.82 4.54 1.82 4.22 4.64 4.22 4.64 1.72 1.82 1.72
                 1.82 1.40 4.96 1.40 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 5.12 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 5.12 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  3.13 2.90 1.46 2.90 1.46 3.68 1.14 3.68 1.14 1.64 1.46 1.64
                 1.46 2.58 3.13 2.58 ;
    END
END buf_8

MACRO buf_64
    CLASS CORE ;
    FOREIGN buf_64 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 29.44 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 5.44  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.47 1.22 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 32.81  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  29.28 4.54 28.96 4.54 28.96 1.72 23.58 1.72 23.58 4.22
                 28.96 4.22 28.96 4.54 23.26 4.54 23.26 1.72 17.98 1.72
                 17.98 4.22 23.26 4.22 23.26 4.54 17.66 4.54 17.66 1.72
                 12.38 1.72 12.38 4.22 17.66 4.22 17.66 4.54 12.06 4.54
                 12.06 1.72 8.47 1.72 8.47 4.22 12.06 4.22 12.06 4.54 6.46 4.54
                 6.46 4.22 8.15 4.22 8.15 1.72 6.46 1.72 6.46 1.40 29.28 1.40 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 29.44 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 29.44 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  7.77 2.90 6.10 2.90 6.10 3.68 5.78 3.68 5.78 1.96 0.48 1.96
                 0.48 3.36 5.78 3.36 5.78 3.68 0.18 3.68 0.18 3.66 0.16 3.66
                 0.16 1.64 6.10 1.64 6.10 2.58 7.77 2.58 ;
    END
END buf_64

MACRO buf_6
    CLASS CORE ;
    FOREIGN buf_6 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.84 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.47 0.68 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.63  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.68 4.30 1.72 4.30 1.72 3.98 3.36 3.98 3.36 1.72 1.73 1.72
                 1.73 1.40 3.68 1.40 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 3.84 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 3.84 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  2.09 2.90 1.36 2.90 1.36 3.68 0.34 3.68 0.34 3.36 1.04 3.36
                 1.04 1.96 0.34 1.96 0.34 1.64 1.36 1.64 1.36 2.58 2.09 2.58 ;
    END
END buf_6

MACRO buf_48
    CLASS CORE ;
    FOREIGN buf_48 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 24.95  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  22.24 4.54 21.92 4.54 21.92 1.72 16.58 1.72 16.58 4.22
                 21.92 4.22 21.92 4.54 16.26 4.54 16.26 1.72 10.98 1.72
                 10.98 4.22 16.26 4.22 16.26 4.54 10.66 4.54 10.66 1.72
                 7.07 1.72 7.07 4.22 10.66 4.22 10.66 4.54 5.06 4.54 5.06 4.22
                 6.75 4.22 6.75 1.72 5.06 1.72 5.06 1.40 22.24 1.40 ;
        END
    END x
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 4.08  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.47 1.22 3.04 ;
        END
    END a
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 22.40 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 22.40 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  6.37 2.90 4.70 2.90 4.70 3.68 4.38 3.68 4.38 1.96 0.48 1.96
                 0.48 3.36 4.38 3.36 4.38 3.68 0.16 3.68 0.16 1.64 4.70 1.64
                 4.70 2.58 6.37 2.58 ;
    END
END buf_48

MACRO buf_4
    CLASS CORE ;
    FOREIGN buf_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.84 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.47 0.78 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.68 4.54 1.82 4.54 1.82 4.22 3.36 4.22 3.36 1.72 1.82 1.72
                 1.82 1.40 3.68 1.40 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 3.84 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 3.84 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  2.82 2.90 1.46 2.90 1.46 4.20 1.14 4.20 1.14 1.34 1.46 1.34
                 1.46 2.58 2.82 2.58 ;
    END
END buf_4

MACRO buf_32
    CLASS CORE ;
    FOREIGN buf_32 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.36 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.72  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.47 1.22 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 17.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  15.20 4.54 14.88 4.54 14.88 1.72 9.58 1.72 9.58 4.22
                 14.88 4.22 14.88 4.54 9.26 4.54 9.26 1.72 5.67 1.72 5.67 4.22
                 9.26 4.22 9.26 4.54 3.66 4.54 3.66 4.22 5.35 4.22 5.35 1.72
                 3.66 1.72 3.66 1.40 15.20 1.40 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 15.36 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 15.36 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.97 2.90 3.30 2.90 3.30 3.68 2.98 3.68 2.98 1.96 0.48 1.96
                 0.48 3.36 2.98 3.36 2.98 3.68 0.16 3.68 0.16 1.64 3.30 1.64
                 3.30 2.58 4.97 2.58 ;
    END
END buf_32

MACRO buf_3
    CLASS CORE ;
    FOREIGN buf_3 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.84 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.47 0.55 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.61  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.68 4.14 1.56 4.14 1.56 3.82 3.36 3.82 3.36 1.65 1.57 1.65
                 1.57 1.33 3.68 1.33 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 3.84 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 3.84 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  1.91 2.90 1.20 2.90 1.20 4.20 0.18 4.20 0.18 3.88 0.88 3.88
                 0.88 1.66 0.18 1.66 0.18 1.34 1.20 1.34 1.20 2.58 1.91 2.58 ;
    END
END buf_3

MACRO buf_24
    CLASS CORE ;
    FOREIGN buf_24 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.16 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.04  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.47 1.46 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 13.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  12.00 4.54 11.68 4.54 11.68 1.72 5.23 1.72 5.23 4.22
                 11.68 4.22 11.68 4.54 3.22 4.54 3.22 4.22 4.91 4.22 4.91 1.72
                 3.22 1.72 3.22 1.40 12.00 1.40 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 12.16 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 12.16 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.53 2.90 2.86 2.90 2.86 3.68 1.13 3.68 1.13 3.36 2.54 3.36
                 2.54 1.96 1.13 1.96 1.13 1.64 2.86 1.64 2.86 2.58 4.53 2.58 ;
    END
END buf_24

MACRO buf_20
    CLASS CORE ;
    FOREIGN buf_20 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.88 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.04  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.47 1.46 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 11.19  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  10.72 4.54 10.40 4.54 10.40 1.72 5.23 1.72 5.23 4.22
                 10.40 4.22 10.40 4.54 3.22 4.54 3.22 4.22 4.91 4.22 4.91 1.72
                 3.22 1.72 3.22 1.40 10.72 1.40 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 10.88 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 10.88 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.53 2.90 2.86 2.90 2.86 3.68 1.13 3.68 1.13 3.36 2.54 3.36
                 2.54 1.96 1.13 1.96 1.13 1.64 2.86 1.64 2.86 2.58 4.53 2.58 ;
    END
END buf_20

MACRO buf_2
    CLASS CORE ;
    FOREIGN buf_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.56 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.78 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  2.40 4.54 1.82 4.54 1.82 4.22 2.08 4.22 2.08 1.54 1.82 1.54
                 1.82 1.22 2.40 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  2.56 0.90 1.28 0.90 1.28 1.72 0.96 1.72 0.96 0.90 0.00 0.90
                 0.00 -0.90 2.56 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  2.56 6.66 0.00 6.66 0.00 4.86 0.98 4.86 0.98 4.34 1.30 4.34
                 1.30 4.86 2.56 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  1.76 3.42 0.48 3.42 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 3.10 1.44 3.10
                 1.44 2.59 1.76 2.59 ;
    END
END buf_2

MACRO buf_16
    CLASS CORE ;
    FOREIGN buf_16 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.96 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.47 1.36 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 9.22  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.30 1.72 8.16 1.72 8.16 4.22 8.30 4.22 8.30 4.54 7.84 4.54
                 7.84 1.72 4.39 1.72 4.39 4.22 7.84 4.22 7.84 4.54 2.38 4.54
                 2.38 4.22 4.07 4.22 4.07 1.72 2.38 1.72 2.38 1.40 8.30 1.40 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 8.96 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 8.96 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  3.69 2.90 2.02 2.90 2.02 3.68 0.29 3.68 0.29 3.36 1.70 3.36
                 1.70 1.96 0.29 1.96 0.29 1.64 2.02 1.64 2.02 2.58 3.69 2.58 ;
    END
END buf_16

MACRO buf_12
    CLASS CORE ;
    FOREIGN buf_12 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.47 1.36 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 7.26  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  6.92 4.54 2.38 4.54 2.38 4.22 6.60 4.22 6.60 3.04 6.56 3.04
                 6.56 2.72 6.60 2.72 6.60 1.72 2.38 1.72 2.38 1.40 6.92 1.40 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 7.68 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 7.68 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  3.69 2.90 2.02 2.90 2.02 3.68 0.29 3.68 0.29 3.36 1.70 3.36
                 1.70 1.96 0.29 1.96 0.29 1.64 2.02 1.64 2.02 2.58 3.69 2.58 ;
    END
END buf_12

MACRO buf_10
    CLASS CORE ;
    FOREIGN buf_10 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.04 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.47 1.36 3.04 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.59  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  5.60 4.54 2.38 4.54 2.38 4.22 5.28 4.22 5.28 1.72 2.38 1.72
                 2.38 1.40 5.60 1.40 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 7.04 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 7.04 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  3.69 2.90 2.02 2.90 2.02 3.68 0.29 3.68 0.29 3.36 1.70 3.36
                 1.70 1.96 0.29 1.96 0.29 1.64 2.02 1.64 2.02 2.58 3.69 2.58 ;
    END
END buf_10

MACRO buf_1
    CLASS CORE ;
    FOREIGN buf_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.56 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.45  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.44 2.41 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  2.40 4.54 1.82 4.54 1.82 4.22 2.08 4.22 2.08 1.54 1.82 1.54
                 1.82 1.22 2.40 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 2.56 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  2.56 6.66 0.00 6.66 0.00 4.86 0.98 4.86 0.98 4.34 1.30 4.34
                 1.30 4.86 2.56 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  1.72 3.55 0.48 3.55 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 3.23 1.72 3.23 ;
    END
END buf_1

MACRO buf_0
    CLASS CORE ;
    FOREIGN buf_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.56 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.45  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.44 2.41 ;
        END
    END a
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.10  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  2.40 4.54 1.82 4.54 1.82 4.22 2.08 4.22 2.08 1.54 1.82 1.54
                 1.82 1.22 2.40 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 2.56 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  2.56 6.66 0.00 6.66 0.00 4.86 0.98 4.86 0.98 4.34 1.30 4.34
                 1.30 4.86 2.56 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  1.72 3.77 0.48 3.77 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 3.45 1.72 3.45 ;
    END
END buf_0

MACRO aoi33_4
    CLASS CORE ;
    FOREIGN aoi33_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.16 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  10.40 2.58 10.72 3.22 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  8.48 2.58 8.80 3.22 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  7.20 2.58 7.52 3.22 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.58 1.12 3.22 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.58 3.04 3.22 ;
        END
    END e
    PIN f
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 2.58 5.60 3.22 ;
        END
    END f
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 7.26  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.46 2.18 4.96 2.18 4.96 3.54 5.36 3.54 5.36 3.86 0.50 3.86
                 0.50 4.50 0.18 4.50 0.18 3.54 4.64 3.54 4.64 2.18 4.34 2.18
                 4.34 1.86 5.74 1.86 5.74 1.22 6.06 1.22 6.06 1.86 7.46 1.86 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 12.16 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  12.16 6.66 0.00 6.66 0.00 4.86 7.12 4.86 7.12 4.18 7.44 4.18
                 7.44 4.86 8.52 4.86 8.52 4.18 8.84 4.18 8.84 4.86 10.60 4.86
                 10.60 4.18 10.92 4.18 10.92 4.86 12.16 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  8.52 1.22 11.62 1.54 ;
        POLYGON  11.62 4.50 11.30 4.50 11.30 3.86 10.22 3.86 10.22 4.50
                 9.90 4.50 9.90 3.86 9.54 3.86 9.54 4.50 9.22 4.50 9.22 3.86
                 8.14 3.86 8.14 4.50 7.82 4.50 7.82 3.86 6.74 3.86 6.74 4.50
                 6.42 4.50 6.42 3.86 6.06 3.86 6.06 4.50 0.88 4.50 0.88 4.18
                 5.74 4.18 5.74 3.54 11.62 3.54 ;
        POLYGON  9.54 2.18 7.82 2.18 7.82 1.54 6.44 1.54 6.44 1.22 8.14 1.22
                 8.14 1.86 9.54 1.86 ;
        POLYGON  5.36 1.54 3.98 1.54 3.98 2.18 2.26 2.18 2.26 1.86 3.66 1.86
                 3.66 1.22 5.36 1.22 ;
        RECT  0.18 1.22 3.28 1.54 ;
    END
END aoi33_4

MACRO aoi33_2
    CLASS CORE ;
    FOREIGN aoi33_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.58 6.88 3.22 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 2.58 5.60 3.22 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.58 4.96 3.22 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.58 0.48 3.22 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.58 1.76 3.22 ;
        END
    END e
    PIN f
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.58 3.68 3.22 ;
        END
    END f
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.76  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.32 3.86 0.50 3.86 0.50 4.50 0.18 4.50 0.18 3.54 4.00 3.54
                 4.00 2.20 3.64 2.20 3.64 1.46 3.96 1.46 3.96 1.88 4.32 1.88 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 7.68 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 6.66 0.00 6.66 0.00 4.86 5.72 4.86 5.72 4.18 6.04 4.18
                 6.04 4.86 6.40 4.86 6.40 4.18 6.72 4.18 6.72 4.86 7.68 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  5.72 1.22 7.42 1.54 ;
        POLYGON  7.42 4.50 7.10 4.50 7.10 3.86 5.34 3.86 5.34 4.50 0.88 4.50
                 0.88 4.18 5.02 4.18 5.02 3.54 7.42 3.54 ;
        RECT  4.34 1.22 5.34 1.54 ;
        RECT  2.26 1.22 3.26 1.54 ;
        RECT  0.18 1.22 1.88 1.54 ;
    END
END aoi33_2

MACRO aoi33_1
    CLASS CORE ;
    FOREIGN aoi33_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.53  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.58 6.88 3.22 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.53  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 2.58 5.60 3.22 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.53  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.58 4.96 3.22 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.53  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.58 0.48 3.22 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.53  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.58 1.76 3.22 ;
        END
    END e
    PIN f
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.53  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.58 3.68 3.22 ;
        END
    END f
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.82  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.96 2.20 3.04 2.20 3.04 3.54 3.26 3.54 3.26 3.86 0.50 3.86
                 0.50 4.50 0.18 4.50 0.18 3.54 2.72 3.54 2.72 1.88 3.96 1.88 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 0.90 6.72 0.90 6.72 1.20 6.40 1.20 6.40 0.90 1.20 0.90
                 1.20 1.20 0.88 1.20 0.88 0.90 0.00 0.90 0.00 -0.90 7.68 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 6.66 0.00 6.66 0.00 4.86 4.32 4.86 4.32 4.78 4.64 4.78
                 4.64 4.86 5.72 4.86 5.72 4.78 6.72 4.78 6.72 4.86 7.68 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  7.42 2.20 5.72 2.20 5.72 1.22 6.04 1.22 6.04 1.88 7.42 1.88 ;
        POLYGON  7.42 4.46 3.96 4.46 3.96 4.50 0.88 4.50 0.88 4.18 3.64 4.18
                 3.64 4.14 7.42 4.14 ;
        RECT  4.34 1.22 5.34 1.54 ;
        RECT  2.26 1.22 3.26 1.54 ;
        POLYGON  1.88 2.20 0.18 2.20 0.18 1.88 1.56 1.88 1.56 1.22 1.88 1.22 ;
    END
END aoi33_1

MACRO aoi32_4
    CLASS CORE ;
    FOREIGN aoi32_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.24 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  8.48 2.54 8.80 3.18 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.54 6.88 3.18 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 2.54 5.60 3.18 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.54 3.68 3.18 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.54 1.12 3.18 ;
        END
    END e
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.29  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  5.38 2.18 4.96 2.18 4.96 3.82 0.50 3.82 0.50 4.50 0.18 4.50
                 0.18 3.50 4.64 3.50 4.64 2.18 2.26 2.18 2.26 1.86 3.66 1.86
                 3.66 1.22 3.98 1.22 3.98 1.86 5.38 1.86 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 10.24 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  10.24 6.66 0.00 6.66 0.00 4.86 6.44 4.86 6.44 4.18 6.76 4.18
                 6.76 4.86 8.52 4.86 8.52 4.18 8.84 4.18 8.84 4.86 10.24 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  6.44 1.22 9.54 1.54 ;
        POLYGON  9.54 4.50 9.22 4.50 9.22 3.82 8.14 3.82 8.14 4.50 7.82 4.50
                 7.82 3.82 7.46 3.82 7.46 4.50 7.14 4.50 7.14 3.82 6.06 3.82
                 6.06 4.50 0.88 4.50 0.88 4.18 5.74 4.18 5.74 3.50 9.54 3.50 ;
        POLYGON  7.46 2.18 5.74 2.18 5.74 1.54 4.36 1.54 4.36 1.22 6.06 1.22
                 6.06 1.86 7.46 1.86 ;
        RECT  0.18 1.22 3.28 1.54 ;
    END
END aoi32_4

MACRO aoi32_2
    CLASS CORE ;
    FOREIGN aoi32_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 2.54 5.60 3.18 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.54 4.32 3.18 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.54 3.68 3.18 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.54 2.40 3.18 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.54 1.12 3.18 ;
        END
    END e
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.77  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.04 3.82 0.50 3.82 0.50 4.50 0.18 4.50 0.18 3.50 2.72 3.50
                 2.72 2.18 2.26 2.18 2.26 1.22 2.58 1.22 2.58 1.86 3.04 1.86 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 6.40 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 6.66 0.00 6.66 0.00 4.86 4.34 4.86 4.34 4.18 5.34 4.18
                 5.34 4.86 6.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  4.34 1.22 6.04 1.54 ;
        POLYGON  6.04 4.50 5.72 4.50 5.72 3.82 3.96 3.82 3.96 4.50 0.88 4.50
                 0.88 4.18 3.64 4.18 3.64 3.50 6.04 3.50 ;
        RECT  2.96 1.22 3.96 1.54 ;
        RECT  0.18 1.22 1.88 1.54 ;
    END
END aoi32_2

MACRO aoi32_1
    CLASS CORE ;
    FOREIGN aoi32_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 2.62 5.60 3.26 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.62 4.32 3.26 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.62 3.68 3.26 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.54 2.40 3.18 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.54 1.12 3.18 ;
        END
    END e
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.99  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.04 3.82 0.18 3.82 0.18 3.50 2.72 3.50 2.72 2.18 2.26 2.18
                 2.26 1.22 2.58 1.22 2.58 1.86 3.04 1.86 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 0.90 5.34 0.90 5.34 1.20 5.02 1.20 5.02 0.90 1.20 0.90
                 1.20 1.20 0.88 1.20 0.88 0.90 0.00 0.90 0.00 -0.90 6.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 6.40 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  6.04 1.96 4.34 1.96 4.34 1.22 4.66 1.22 4.66 1.64 6.04 1.64 ;
        RECT  0.88 4.18 6.04 4.50 ;
        RECT  2.96 1.22 3.96 1.54 ;
        POLYGON  1.88 1.96 0.18 1.96 0.18 1.64 1.56 1.64 1.56 1.22 1.88 1.22 ;
    END
END aoi32_1

MACRO aoi31_4
    CLASS CORE ;
    FOREIGN aoi31_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.62 6.88 3.26 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.62 4.96 3.26 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.62 3.04 3.26 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.62 1.12 3.26 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 7.31  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.46 4.54 7.14 4.54 7.14 3.90 0.16 3.90 0.16 1.22 1.90 1.22
                 1.90 1.86 3.30 1.86 3.30 2.18 1.58 2.18 1.58 1.54 0.48 1.54
                 0.48 3.58 7.46 3.58 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 7.68 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 7.68 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  7.46 1.54 5.38 1.54 5.38 2.18 3.66 2.18 3.66 1.86 5.06 1.86
                 5.06 1.22 7.46 1.22 ;
        RECT  0.18 4.22 6.76 4.54 ;
        RECT  2.28 1.22 4.68 1.54 ;
    END
END aoi31_4

MACRO aoi31_2
    CLASS CORE ;
    FOREIGN aoi31_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.08 4.32 2.72 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.08 3.04 2.72 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.08 2.40 2.72 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.72 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.95  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.52 3.90 0.16 3.90 0.16 1.22 1.44 1.22 1.44 1.54 0.48 1.54
                 0.48 3.58 3.52 3.58 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 5.12 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 6.66 0.00 6.66 0.00 4.86 0.42 4.86 0.42 4.22 0.74 4.22
                 0.74 4.86 5.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  3.20 1.22 4.90 1.54 ;
        POLYGON  4.22 4.54 1.12 4.54 1.12 4.22 3.90 4.22 3.90 3.58 4.22 3.58 ;
        RECT  1.82 1.22 2.82 1.54 ;
    END
END aoi31_2

MACRO aoi31_1
    CLASS CORE ;
    FOREIGN aoi31_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.08 4.32 2.72 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.08 3.04 2.72 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.08 2.40 2.72 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.72 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.12  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.52 3.90 0.16 3.90 0.16 1.22 1.44 1.22 1.44 1.54 0.48 1.54
                 0.48 3.58 3.52 3.58 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 5.12 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 6.66 0.00 6.66 0.00 4.86 0.42 4.86 0.42 4.22 0.74 4.22
                 0.74 4.86 5.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  3.20 1.22 4.90 1.54 ;
        RECT  1.12 4.22 4.22 4.54 ;
        RECT  1.82 1.22 2.82 1.54 ;
    END
END aoi31_1

MACRO aoi22_4
    CLASS CORE ;
    FOREIGN aoi22_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.62 1.12 3.26 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.62 3.04 3.26 ;
        END
    END b
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.92 2.62 6.24 3.26 ;
        END
    END d
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.62 4.96 3.26 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.29  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  6.80 4.54 6.48 4.54 6.48 3.90 3.36 3.90 3.36 2.18 2.26 2.18
                 2.26 1.86 3.66 1.86 3.66 1.22 3.98 1.22 3.98 1.86 5.38 1.86
                 5.38 2.18 3.68 2.18 3.68 3.58 6.80 3.58 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 7.68 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 7.68 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  4.36 1.22 7.46 1.54 ;
        POLYGON  6.10 4.54 1.58 4.54 1.58 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 3.58 1.90 3.58 1.90 4.22 6.10 4.22 ;
        RECT  0.18 1.22 3.28 1.54 ;
    END
END aoi22_4

MACRO aoi22_2
    CLASS CORE ;
    FOREIGN aoi22_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.62 1.12 3.26 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.62 1.76 3.26 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.62 3.04 3.26 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.62 4.32 3.26 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.97  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.52 3.90 2.08 3.90 2.08 1.98 2.26 1.98 2.26 1.22 2.58 1.22
                 2.58 2.30 2.40 2.30 2.40 3.58 3.52 3.58 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 0.90 4.66 0.90 4.66 1.54 4.34 1.54 4.34 0.90 0.00 0.90
                 0.00 -0.90 5.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 6.66 0.00 6.66 0.00 4.86 0.42 4.86 0.42 3.66 0.74 3.66
                 0.74 4.86 5.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.22 4.54 1.12 4.54 1.12 3.66 1.44 3.66 1.44 4.22 3.90 4.22
                 3.90 3.66 4.22 3.66 ;
        RECT  2.96 1.22 3.96 1.54 ;
        RECT  0.18 1.22 1.88 1.54 ;
    END
END aoi22_2

MACRO aoi22_1
    CLASS CORE ;
    FOREIGN aoi22_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.48 2.72 1.12 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.72 2.08 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.72 3.04 3.04 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.72 4.64 3.04 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.41  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.68 3.90 3.20 3.90 3.20 3.58 3.36 3.58 3.36 2.40 2.26 2.40
                 2.26 1.74 2.58 1.74 2.58 2.08 3.68 2.08 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 0.90 4.66 0.90 4.66 1.76 4.34 1.76 4.34 0.90 1.20 0.90
                 1.20 1.30 0.88 1.30 0.88 0.90 0.00 0.90 0.00 -0.90 5.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 6.66 0.00 6.66 0.00 4.86 0.42 4.86 0.42 4.52 0.74 4.52
                 0.74 4.86 1.82 4.86 1.82 4.52 2.14 4.52 2.14 4.86 5.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.22 4.54 2.50 4.54 2.50 4.20 1.12 4.20 1.12 3.88 2.82 3.88
                 2.82 4.22 4.22 4.22 ;
        RECT  2.96 1.44 3.96 1.76 ;
        POLYGON  1.88 2.08 0.18 2.08 0.18 1.44 0.50 1.44 0.50 1.76 1.56 1.76
                 1.56 1.44 1.88 1.44 ;
    END
END aoi22_1

MACRO aoi222_4
    CLASS CORE ;
    FOREIGN aoi222_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.52 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  7.84 2.50 8.16 3.14 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.50 4.96 3.14 ;
        END
    END c
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  9.76 2.50 10.08 3.14 ;
        END
    END a
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.50 6.88 3.14 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.50 3.04 3.14 ;
        END
    END e
    PIN f
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.50 1.12 3.14 ;
        END
    END f
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.86 2.18 1.76 2.18 1.76 3.54 3.30 3.54 3.30 3.86 0.50 3.86
                 0.50 4.54 0.18 4.54 0.18 3.54 1.44 3.54 1.44 2.18 0.18 2.18
                 0.18 1.22 0.50 1.22 0.50 1.86 7.14 1.86 7.14 1.22 7.46 1.22
                 7.46 1.86 8.86 1.86 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  11.52 0.90 10.24 0.90 10.24 1.54 9.92 1.54 9.92 0.90 3.98 0.90
                 3.98 1.54 3.66 1.54 3.66 0.90 0.00 0.90 0.00 -0.90 11.52 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  11.52 6.66 0.00 6.66 0.00 4.86 8.52 4.86 8.52 4.22 8.84 4.22
                 8.84 4.86 9.92 4.86 9.92 4.22 10.24 4.22 10.24 4.86 11.52 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  10.94 2.18 9.22 2.18 9.22 1.54 7.84 1.54 7.84 1.22 9.54 1.22
                 9.54 1.86 10.62 1.86 10.62 1.22 10.94 1.22 ;
        POLYGON  10.94 4.54 10.62 4.54 10.62 3.86 9.54 3.86 9.54 4.54 9.22 4.54
                 9.22 3.86 8.14 3.86 8.14 4.54 7.82 4.54 7.82 3.86 3.66 3.86
                 3.66 3.54 10.94 3.54 ;
        RECT  0.88 4.22 7.46 4.54 ;
        RECT  4.36 1.22 6.76 1.54 ;
        RECT  0.88 1.22 3.28 1.54 ;
    END
END aoi222_4

MACRO aoi222_2
    CLASS CORE ;
    FOREIGN aoi222_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.88 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.08  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  9.12 2.50 9.44 3.14 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.08  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  7.84 2.50 8.16 3.14 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.08  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.50 4.96 3.14 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.08  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.92 2.50 6.24 3.14 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.08  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.50 2.40 3.14 ;
        END
    END e
    PIN f
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.08  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.50 1.12 3.14 ;
        END
    END f
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.17  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.46 2.18 3.04 2.18 3.04 3.54 3.30 3.54 3.30 3.86 0.18 3.86
                 0.18 3.54 2.72 3.54 2.72 2.18 0.18 2.18 0.18 1.22 0.50 1.22
                 0.50 1.86 5.76 1.86 5.76 1.22 6.08 1.22 6.08 1.86 7.14 1.86
                 7.14 1.22 7.46 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  10.88 0.90 8.86 0.90 8.86 1.54 8.54 1.54 8.54 0.90 3.98 0.90
                 3.98 1.54 3.66 1.54 3.66 0.90 2.60 0.90 2.60 1.54 2.28 1.54
                 2.28 0.90 0.00 0.90 0.00 -0.90 10.88 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  10.88 6.66 0.00 6.66 0.00 4.86 7.84 4.86 7.84 4.22 8.16 4.22
                 8.16 4.86 9.24 4.86 9.24 4.22 9.56 4.22 9.56 4.86 10.88 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  10.26 4.54 9.94 4.54 9.94 3.86 8.86 3.86 8.86 4.54 8.54 4.54
                 8.54 3.86 7.46 3.86 7.46 4.54 7.14 4.54 7.14 3.86 3.66 3.86
                 3.66 3.54 10.26 3.54 ;
        POLYGON  9.56 2.18 7.84 2.18 7.84 1.22 8.16 1.22 8.16 1.86 9.24 1.86
                 9.24 1.22 9.56 1.22 ;
        RECT  0.88 4.22 6.08 4.54 ;
        RECT  4.36 1.22 5.38 1.54 ;
        RECT  0.88 1.22 1.90 1.54 ;
    END
END aoi222_2

MACRO aoi222_1
    CLASS CORE ;
    FOREIGN aoi222_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.04 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.92 2.72 6.56 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.72 5.28 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.36 3.04 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.68 2.72 4.32 3.04 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.72 2.08 3.04 ;
        END
    END e
    PIN f
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.48 3.36 ;
        END
    END f
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.16  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.66 2.18 1.12 2.18 1.12 3.54 1.52 3.54 1.52 3.86 0.80 3.86
                 0.80 2.18 0.18 2.18 0.18 1.22 0.50 1.22 0.50 1.86 4.34 1.86
                 4.34 1.22 4.66 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  7.04 0.90 6.04 0.90 6.04 1.54 5.72 1.54 5.72 0.90 2.58 0.90
                 2.58 1.54 2.26 1.54 2.26 0.90 0.00 0.90 0.00 -0.90 7.04 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.04 6.66 0.00 6.66 0.00 4.86 5.60 4.86 5.60 4.22 5.92 4.22
                 5.92 4.86 7.04 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  6.74 2.18 5.04 2.18 5.04 1.22 5.36 1.22 5.36 1.86 6.42 1.86
                 6.42 1.22 6.74 1.22 ;
        POLYGON  6.62 4.54 6.30 4.54 6.30 3.86 5.22 3.86 5.22 4.54 4.90 4.54
                 4.90 3.86 3.44 3.86 3.44 3.54 6.62 3.54 ;
        POLYGON  4.54 4.54 0.42 4.54 0.42 4.22 2.66 4.22 2.66 3.54 2.98 3.54
                 2.98 4.22 4.54 4.22 ;
        RECT  2.96 1.22 3.96 1.54 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END aoi222_1

MACRO aoi221_4
    CLASS CORE ;
    FOREIGN aoi221_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.24 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  8.48 2.50 8.80 3.14 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.50 6.88 3.14 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.50 3.04 3.14 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.50 0.48 3.14 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 2.50 5.60 3.14 ;
        END
    END e
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.46 2.18 1.76 2.18 1.76 3.54 3.30 3.54 3.30 3.86 0.50 3.86
                 0.50 4.54 0.18 4.54 0.18 3.54 1.44 3.54 1.44 2.18 0.18 2.18
                 0.18 1.22 0.50 1.22 0.50 1.86 4.34 1.86 4.34 1.22 4.66 1.22
                 4.66 1.86 5.74 1.86 5.74 1.22 6.06 1.22 6.06 1.86 7.46 1.86 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  10.24 0.90 5.36 0.90 5.36 1.54 5.04 1.54 5.04 0.90 3.98 0.90
                 3.98 1.54 3.66 1.54 3.66 0.90 0.00 0.90 0.00 -0.90 10.24 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  10.24 6.66 0.00 6.66 0.00 4.86 6.44 4.86 6.44 4.22 6.76 4.22
                 6.76 4.86 8.52 4.86 8.52 4.22 8.84 4.22 8.84 4.86 10.24 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  6.44 1.22 9.54 1.54 ;
        POLYGON  9.54 4.54 9.22 4.54 9.22 3.86 8.14 3.86 8.14 4.54 7.82 4.54
                 7.82 3.86 7.46 3.86 7.46 4.54 7.14 4.54 7.14 3.86 6.06 3.86
                 6.06 4.54 4.36 4.54 4.36 4.22 5.74 4.22 5.74 3.54 9.54 3.54 ;
        POLYGON  5.38 3.86 3.98 3.86 3.98 4.54 0.88 4.54 0.88 4.22 3.66 4.22
                 3.66 3.54 5.38 3.54 ;
        RECT  0.88 1.22 3.28 1.54 ;
    END
END aoi221_4

MACRO aoi221_2
    CLASS CORE ;
    FOREIGN aoi221_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.76 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.50 4.96 3.14 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.50 3.68 3.14 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.50 1.76 3.14 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.50 0.48 3.14 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.50 3.04 3.14 ;
        END
    END e
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.45  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.28 2.18 2.40 2.18 2.40 3.86 0.50 3.86 0.50 4.54 0.18 4.54
                 0.18 3.54 2.08 3.54 2.08 2.18 0.18 2.18 0.18 1.22 0.50 1.22
                 0.50 1.86 2.96 1.86 2.96 1.22 3.28 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  5.76 0.90 2.58 0.90 2.58 1.54 2.26 1.54 2.26 0.90 0.00 0.90
                 0.00 -0.90 5.76 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.76 6.66 0.00 6.66 0.00 4.86 4.34 4.86 4.34 4.22 4.66 4.22
                 4.66 4.86 5.76 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  3.66 1.22 5.36 1.54 ;
        POLYGON  5.36 4.54 5.04 4.54 5.04 3.86 3.96 3.86 3.96 4.54 2.96 4.54
                 2.96 3.54 5.36 3.54 ;
        RECT  0.88 4.22 2.58 4.54 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END aoi221_2

MACRO aoi221_1
    CLASS CORE ;
    FOREIGN aoi221_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.76 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.50 4.96 3.14 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.50 3.68 3.14 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.50 1.76 3.14 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.50 0.48 3.14 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.50 3.04 3.14 ;
        END
    END e
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.48  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.28 2.18 2.40 2.18 2.40 3.86 0.18 3.86 0.18 3.54 2.08 3.54
                 2.08 2.18 0.18 2.18 0.18 1.22 0.50 1.22 0.50 1.86 2.96 1.86
                 2.96 1.22 3.28 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  5.76 0.90 4.66 0.90 4.66 1.20 4.34 1.20 4.34 0.90 2.58 0.90
                 2.58 1.54 2.26 1.54 2.26 0.90 0.00 0.90 0.00 -0.90 5.76 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.76 6.66 0.00 6.66 0.00 4.86 4.34 4.86 4.34 4.78 4.66 4.78
                 4.66 4.86 5.76 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  5.36 1.84 3.66 1.84 3.66 1.22 3.98 1.22 3.98 1.52 5.04 1.52
                 5.04 1.22 5.36 1.22 ;
        POLYGON  5.36 4.54 5.04 4.54 5.04 4.46 3.96 4.46 3.96 4.54 2.96 4.54
                 2.96 4.22 3.64 4.22 3.64 4.14 5.36 4.14 ;
        RECT  0.88 4.22 2.58 4.54 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END aoi221_1

MACRO aoi21_4
    CLASS CORE ;
    FOREIGN aoi21_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.76 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.08 4.96 2.72 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.62 3.36 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.72 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.34  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  5.38 4.54 5.06 4.54 5.06 3.90 0.16 3.90 0.16 1.22 3.30 1.22
                 3.30 1.54 0.48 1.54 0.48 3.58 5.38 3.58 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 5.76 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 5.76 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  5.38 1.54 3.98 1.54 3.98 2.18 2.16 2.18 2.16 1.86 3.66 1.86
                 3.66 1.22 5.38 1.22 ;
        RECT  0.18 4.22 4.68 4.54 ;
    END
END aoi21_4

MACRO aoi21_2
    CLASS CORE ;
    FOREIGN aoi21_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.84 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.08 3.04 2.72 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.08 2.40 2.72 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.72 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.77  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.52 4.32 3.20 4.32 3.20 3.90 0.16 3.90 0.16 1.22 1.44 1.22
                 1.44 1.54 0.48 1.54 0.48 3.58 3.52 3.58 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 3.84 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  3.84 6.66 0.00 6.66 0.00 4.86 0.42 4.86 0.42 4.22 0.74 4.22
                 0.74 4.86 3.84 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  1.82 1.22 3.52 1.54 ;
        RECT  1.12 4.22 2.82 4.54 ;
    END
END aoi21_2

MACRO aoi21_1
    CLASS CORE ;
    FOREIGN aoi21_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.84 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.08 3.04 2.72 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.08 2.40 2.72 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.72 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.99  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.52 4.32 3.20 4.32 3.20 3.90 0.16 3.90 0.16 1.22 1.44 1.22
                 1.44 1.54 0.48 1.54 0.48 3.58 3.52 3.58 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 3.84 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  3.84 6.66 0.00 6.66 0.00 4.86 0.42 4.86 0.42 4.22 0.74 4.22
                 0.74 4.86 3.84 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  1.82 1.22 3.52 1.54 ;
        RECT  1.12 4.22 2.82 4.54 ;
    END
END aoi21_1

MACRO aoi211_4
    CLASS CORE ;
    FOREIGN aoi211_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.50 3.04 3.24 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.50 1.12 3.24 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.50 6.88 3.24 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.50 4.96 3.24 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.65  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.46 2.18 5.74 2.18 5.74 1.54 4.68 1.54 4.68 2.18 1.76 2.18
                 1.76 3.58 3.30 3.58 3.30 3.90 0.50 3.90 0.50 4.54 0.18 4.54
                 0.18 3.58 1.44 3.58 1.44 2.18 0.18 2.18 0.18 1.22 0.50 1.22
                 0.50 1.86 4.36 1.86 4.36 1.22 6.06 1.22 6.06 1.86 7.14 1.86
                 7.14 1.22 7.46 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 0.90 6.76 0.90 6.76 1.54 6.44 1.54 6.44 0.90 3.98 0.90
                 3.98 1.54 3.66 1.54 3.66 0.90 0.00 0.90 0.00 -0.90 7.68 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 6.66 0.00 6.66 0.00 4.86 6.44 4.86 6.44 4.22 6.76 4.22
                 6.76 4.86 7.68 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  7.46 4.54 7.14 4.54 7.14 3.90 6.06 3.90 6.06 4.54 4.36 4.54
                 4.36 4.22 5.74 4.22 5.74 3.58 7.46 3.58 ;
        POLYGON  5.38 3.90 3.98 3.90 3.98 4.54 0.88 4.54 0.88 4.22 3.66 4.22
                 3.66 3.58 5.38 3.58 ;
        RECT  0.88 1.22 3.28 1.54 ;
    END
END aoi211_4

MACRO aoi211_2
    CLASS CORE ;
    FOREIGN aoi211_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.50 1.76 3.24 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.50 0.48 3.24 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.50 4.32 3.24 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.50 3.04 3.24 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.00  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.96 1.54 3.28 1.54 3.28 2.18 1.12 2.18 1.12 3.58 1.90 3.58
                 1.90 3.90 0.50 3.90 0.50 4.54 0.18 4.54 0.18 3.58 0.80 3.58
                 0.80 2.18 0.18 2.18 0.18 1.22 0.50 1.22 0.50 1.86 2.96 1.86
                 2.96 1.22 3.96 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 0.90 4.66 0.90 4.66 1.54 4.34 1.54 4.34 0.90 2.58 0.90
                 2.58 1.54 2.26 1.54 2.26 0.90 0.00 0.90 0.00 -0.90 5.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 6.66 0.00 6.66 0.00 4.86 4.34 4.86 4.34 3.58 4.66 3.58
                 4.66 4.86 5.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  2.96 3.58 3.96 4.54 ;
        POLYGON  2.58 4.54 0.88 4.54 0.88 4.22 2.26 4.22 2.26 3.58 2.58 3.58 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END aoi211_2

MACRO aoi211_1
    CLASS CORE ;
    FOREIGN aoi211_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.50 1.76 3.24 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.50 0.48 3.24 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.50 4.32 3.24 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.50 3.04 3.24 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.89  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.96 1.54 3.28 1.54 3.28 2.18 1.12 2.18 1.12 3.58 1.90 3.58
                 1.90 3.90 0.50 3.90 0.50 4.54 0.18 4.54 0.18 3.58 0.80 3.58
                 0.80 2.18 0.18 2.18 0.18 1.22 0.50 1.22 0.50 1.86 2.96 1.86
                 2.96 1.22 3.96 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 0.90 4.66 0.90 4.66 1.54 4.34 1.54 4.34 0.90 2.58 0.90
                 2.58 1.54 2.26 1.54 2.26 0.90 0.00 0.90 0.00 -0.90 5.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 6.66 0.00 6.66 0.00 4.86 4.34 4.86 4.34 4.22 4.66 4.22
                 4.66 4.86 5.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  2.96 4.22 3.96 4.54 ;
        RECT  0.88 4.22 2.58 4.54 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END aoi211_1

MACRO ao33_4
    CLASS CORE ;
    FOREIGN ao33_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.96 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  7.84 2.08 8.16 2.72 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.08 6.88 2.72 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 2.08 5.60 2.72 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.50 1.86 3.04 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.50 3.04 3.14 ;
        END
    END e
    PIN f
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.50 4.32 3.14 ;
        END
    END f
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  0.52 1.54 0.48 1.54 0.48 4.22 0.52 4.22 0.52 4.54 0.16 4.54
                 0.16 1.22 0.52 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.96 0.90 1.34 0.90 1.34 1.54 1.02 1.54 1.02 0.90 0.00 0.90
                 0.00 -0.90 8.96 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  8.96 6.66 0.00 6.66 0.00 4.86 0.90 4.86 0.90 4.22 1.22 4.22
                 1.22 4.86 5.28 4.86 5.28 4.18 5.60 4.18 5.60 4.86 6.68 4.86
                 6.68 4.18 7.64 4.18 7.64 4.86 8.96 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  6.68 1.22 8.38 1.54 ;
        POLYGON  8.38 4.50 8.06 4.50 8.06 3.86 6.30 3.86 6.30 4.50 5.98 4.50
                 5.98 3.86 4.92 3.86 4.92 4.50 2.41 4.50 2.41 4.18 4.60 4.18
                 4.60 3.54 8.38 3.54 ;
        RECT  5.30 1.22 6.30 1.54 ;
        POLYGON  4.92 2.18 1.12 2.18 1.12 3.54 4.18 3.54 4.18 3.86 1.90 3.86
                 1.90 4.50 1.58 4.50 1.58 3.86 0.80 3.86 0.80 1.86 4.60 1.86
                 4.60 1.46 4.92 1.46 ;
        RECT  3.22 1.22 4.22 1.54 ;
        RECT  1.84 1.22 2.84 1.54 ;
    END
END ao33_4

MACRO ao33_2
    CLASS CORE ;
    FOREIGN ao33_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.96 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  7.84 2.08 8.16 2.72 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.08 6.88 2.72 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 2.08 5.60 2.72 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.50 1.76 3.14 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.50 3.04 3.14 ;
        END
    END e
    PIN f
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.50 4.32 3.14 ;
        END
    END f
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  0.52 1.54 0.48 1.54 0.48 4.22 0.52 4.22 0.52 4.54 0.16 4.54
                 0.16 1.22 0.52 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 8.96 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  8.96 6.66 0.00 6.66 0.00 4.86 5.28 4.86 5.28 4.18 5.60 4.18
                 5.60 4.86 6.68 4.86 6.68 4.18 7.64 4.18 7.64 4.86 8.96 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  6.68 1.22 8.38 1.54 ;
        POLYGON  8.38 4.50 8.06 4.50 8.06 3.86 6.30 3.86 6.30 4.50 5.98 4.50
                 5.98 3.86 4.92 3.86 4.92 4.50 2.41 4.50 2.41 4.18 4.60 4.18
                 4.60 3.54 8.38 3.54 ;
        RECT  5.30 1.22 6.30 1.54 ;
        POLYGON  4.92 2.18 1.12 2.18 1.12 3.54 4.18 3.54 4.18 3.86 0.80 3.86
                 0.80 1.86 4.60 1.86 4.60 1.46 4.92 1.46 ;
        RECT  3.22 1.22 4.22 1.54 ;
        RECT  1.84 1.22 2.84 1.54 ;
    END
END ao33_2

MACRO ao33_1
    CLASS CORE ;
    FOREIGN ao33_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.96 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.53  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  7.20 2.72 7.84 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.53  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.57 6.88 3.21 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.53  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.96 2.72 5.60 3.04 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.53  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.72 2.08 3.04 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.53  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.72 3.04 3.04 ;
        END
    END e
    PIN f
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.53  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.68 2.72 4.42 3.12 ;
        END
    END f
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  0.52 1.54 0.48 1.54 0.48 4.22 0.52 4.22 0.52 4.54 0.16 4.54
                 0.16 1.22 0.52 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 8.96 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  8.96 6.66 0.00 6.66 0.00 4.86 0.90 4.86 0.90 4.82 1.22 4.82
                 1.22 4.86 5.28 4.86 5.28 4.82 5.60 4.82 5.60 4.86 6.92 4.86
                 6.92 4.82 7.24 4.82 7.24 4.86 8.96 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  6.68 1.22 8.38 1.54 ;
        RECT  2.41 4.18 8.38 4.50 ;
        RECT  5.30 1.22 6.30 1.54 ;
        POLYGON  4.92 2.18 1.12 2.18 1.12 3.54 3.87 3.54 3.87 3.86 0.80 3.86
                 0.80 1.86 4.60 1.86 4.60 1.46 4.92 1.46 ;
        RECT  3.22 1.22 4.22 1.54 ;
        RECT  1.84 1.22 2.84 1.54 ;
    END
END ao33_1

MACRO ao32_4
    CLASS CORE ;
    FOREIGN ao32_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.04 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.92 2.08 6.24 2.72 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.08 4.96 2.72 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.08 4.32 2.72 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.50 3.04 3.14 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.60 1.86 3.10 ;
        END
    END e
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  0.52 1.54 0.48 1.54 0.48 4.22 0.52 4.22 0.52 4.54 0.16 4.54
                 0.16 1.22 0.52 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  7.04 0.90 1.25 0.90 1.25 1.54 0.93 1.54 0.93 0.90 0.00 0.90
                 0.00 -0.90 7.04 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.04 6.66 0.00 6.66 0.00 4.86 0.90 4.86 0.90 4.18 1.22 4.18
                 1.22 4.86 3.72 4.86 3.72 4.18 4.04 4.18 4.04 4.86 5.12 4.86
                 5.12 4.18 6.08 4.18 6.08 4.86 7.04 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  5.12 1.22 6.82 1.54 ;
        POLYGON  6.82 4.50 6.50 4.50 6.50 3.86 4.74 3.86 4.74 4.50 4.42 4.50
                 4.42 3.86 3.36 3.86 3.36 4.50 1.58 4.50 1.58 4.18 3.04 4.18
                 3.04 3.54 6.82 3.54 ;
        RECT  3.74 1.22 4.74 1.54 ;
        POLYGON  3.36 2.18 1.12 2.18 1.12 3.54 2.63 3.54 2.63 3.86 0.80 3.86
                 0.80 1.86 3.04 1.86 3.04 1.46 3.36 1.46 ;
        RECT  1.66 1.22 2.66 1.54 ;
    END
END ao32_4

MACRO ao32_2
    CLASS CORE ;
    FOREIGN ao32_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  6.56 2.08 6.88 2.72 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 2.08 5.60 2.72 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.08 4.32 2.72 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.50 3.04 3.14 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.60 1.86 3.10 ;
        END
    END e
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  0.52 1.54 0.48 1.54 0.48 4.22 0.52 4.22 0.52 4.54 0.16 4.54
                 0.16 1.22 0.52 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 7.68 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 6.66 0.00 6.66 0.00 4.86 0.90 4.86 0.90 4.22 1.22 4.22
                 1.22 4.86 3.90 4.86 3.90 4.18 4.22 4.18 4.22 4.86 5.30 4.86
                 5.30 4.18 6.26 4.18 6.26 4.86 7.68 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  5.30 1.22 7.00 1.54 ;
        POLYGON  7.00 4.54 6.68 4.54 6.68 3.86 4.92 3.86 4.92 4.54 4.60 4.54
                 4.60 3.86 3.54 3.86 3.54 4.50 1.58 4.50 1.58 4.18 3.22 4.18
                 3.22 3.54 7.00 3.54 ;
        RECT  3.92 1.22 4.92 1.54 ;
        POLYGON  3.54 2.18 1.12 2.18 1.12 3.54 2.60 3.54 2.60 3.86 0.80 3.86
                 0.80 1.86 3.22 1.86 3.22 1.46 3.54 1.46 ;
        RECT  1.84 1.22 2.84 1.54 ;
    END
END ao32_2

MACRO ao32_1
    CLASS CORE ;
    FOREIGN ao32_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.04 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.60 2.72 6.24 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.32 2.72 4.96 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.72 4.00 3.04 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.72 3.04 3.04 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.72 2.08 3.04 ;
        END
    END e
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  0.52 1.54 0.48 1.54 0.48 4.22 0.52 4.22 0.52 4.54 0.16 4.54
                 0.16 1.22 0.52 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  7.04 0.90 6.06 0.90 6.06 1.08 5.74 1.08 5.74 0.90 1.22 0.90
                 1.22 1.08 0.90 1.08 0.90 0.90 0.00 0.90 0.00 -0.90 7.04 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.04 6.66 0.00 6.66 0.00 4.86 0.90 4.86 0.90 4.82 1.22 4.82
                 1.22 4.86 3.66 4.86 3.66 4.82 3.98 4.82 3.98 4.86 5.30 4.86
                 5.30 4.82 5.62 4.82 5.62 4.86 7.04 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  6.76 1.72 5.06 1.72 5.06 1.22 5.38 1.22 5.38 1.40 6.44 1.40
                 6.44 1.22 6.76 1.22 ;
        RECT  1.58 4.18 6.76 4.50 ;
        RECT  3.68 1.22 4.68 1.54 ;
        POLYGON  3.30 2.18 1.12 2.18 1.12 3.54 2.60 3.54 2.60 3.86 0.80 3.86
                 0.80 1.86 2.98 1.86 2.98 1.46 3.30 1.46 ;
        RECT  1.60 1.22 2.60 1.54 ;
    END
END ao32_1

MACRO ao31_4
    CLASS CORE ;
    FOREIGN ao31_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.53  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.62 4.96 3.26 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.53  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.57 3.68 3.21 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.53  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.57 3.04 3.21 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.72 1.86 3.26 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  0.52 1.54 0.48 1.54 0.48 4.22 0.52 4.22 0.52 4.54 0.16 4.54
                 0.16 1.22 0.52 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 6.40 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 6.40 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  1.84 4.22 4.94 4.54 ;
        RECT  3.92 1.46 4.92 1.78 ;
        POLYGON  4.24 3.90 0.80 3.90 0.80 1.98 1.84 1.98 1.84 1.22 2.16 1.22
                 2.16 2.30 1.12 2.30 1.12 3.58 4.24 3.58 ;
        RECT  2.54 1.46 3.54 1.78 ;
    END
END ao31_4

MACRO ao31_2
    CLASS CORE ;
    FOREIGN ao31_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.76 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.53  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.62 4.96 3.26 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.53  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.57 3.70 3.21 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.53  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.57 3.04 3.21 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.72 1.86 3.26 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  0.52 1.54 0.48 1.54 0.48 4.22 0.52 4.22 0.52 4.54 0.16 4.54
                 0.16 1.22 0.52 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 5.76 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 5.76 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  3.68 1.46 5.38 1.78 ;
        RECT  1.84 4.22 4.94 4.54 ;
        POLYGON  4.24 3.90 0.80 3.90 0.80 1.98 1.60 1.98 1.60 1.22 1.92 1.22
                 1.92 2.30 1.12 2.30 1.12 3.58 4.24 3.58 ;
        RECT  2.30 1.46 3.30 1.78 ;
    END
END ao31_2

MACRO ao31_1
    CLASS CORE ;
    FOREIGN ao31_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.76 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.62 4.96 3.26 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.57 3.70 3.21 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.57 3.04 3.21 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.72 1.86 3.26 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  0.52 1.54 0.48 1.54 0.48 4.22 0.52 4.22 0.52 4.54 0.16 4.54
                 0.16 1.22 0.52 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 5.76 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 5.76 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  3.68 1.22 5.38 1.54 ;
        RECT  1.84 4.22 4.94 4.54 ;
        POLYGON  4.24 3.90 0.80 3.90 0.80 1.98 1.60 1.98 1.60 1.22 1.92 1.22
                 1.92 2.30 1.12 2.30 1.12 3.58 4.24 3.58 ;
        RECT  2.30 1.22 3.30 1.54 ;
    END
END ao31_1

MACRO ao22_4
    CLASS CORE ;
    FOREIGN ao22_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.48 2.72 1.12 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.40 1.76 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.72 3.04 3.04 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.40 4.32 3.04 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 1.77 5.60 4.54 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 0.90 4.76 0.90 4.76 1.76 4.44 1.76 4.44 0.90 1.20 0.90
                 1.20 1.30 0.88 1.30 0.88 0.90 0.00 0.90 0.00 -0.90 6.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 6.66 0.00 6.66 0.00 4.86 0.42 4.86 0.42 4.22 0.74 4.22
                 0.74 4.86 1.82 4.86 1.82 4.22 2.14 4.22 2.14 4.86 4.58 4.86
                 4.58 4.22 4.90 4.22 4.90 4.86 6.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.96 3.90 3.20 3.90 3.20 3.58 3.36 3.58 3.36 2.40 2.26 2.40
                 2.26 1.74 2.58 1.74 2.58 2.08 3.68 2.08 3.68 3.58 4.64 3.58
                 4.64 2.62 4.96 2.62 ;
        POLYGON  4.22 4.54 2.50 4.54 2.50 3.90 1.44 3.90 1.44 4.54 1.12 4.54
                 1.12 3.58 2.82 3.58 2.82 4.22 4.22 4.22 ;
        RECT  2.96 1.44 3.96 1.76 ;
        POLYGON  1.88 2.08 0.18 2.08 0.18 1.44 0.50 1.44 0.50 1.76 1.56 1.76
                 1.56 1.44 1.88 1.44 ;
    END
END ao22_4

MACRO ao22_2
    CLASS CORE ;
    FOREIGN ao22_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.76 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.48 2.72 1.12 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.40 1.76 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.72 3.04 3.04 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.40 4.32 3.04 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  5.60 4.54 5.26 4.54 5.26 4.22 5.28 4.22 5.28 2.09 5.26 2.09
                 5.26 1.77 5.60 1.77 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  5.76 0.90 4.84 0.90 4.84 1.76 4.52 1.76 4.52 0.90 1.20 0.90
                 1.20 1.30 0.88 1.30 0.88 0.90 0.00 0.90 0.00 -0.90 5.76 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.76 6.66 0.00 6.66 0.00 4.86 1.10 4.86 1.10 4.22 1.42 4.22
                 1.42 4.86 4.56 4.86 4.56 4.22 4.88 4.22 4.88 4.86 5.76 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.96 3.90 3.18 3.90 3.18 3.58 3.36 3.58 3.36 2.40 2.26 2.40
                 2.26 1.74 2.58 1.74 2.58 2.08 3.68 2.08 3.68 3.58 4.64 3.58
                 4.64 3.08 4.96 3.08 ;
        POLYGON  4.20 4.54 2.48 4.54 2.48 3.90 2.12 3.90 2.12 4.54 1.80 4.54
                 1.80 3.90 0.72 3.90 0.72 4.54 0.40 4.54 0.40 3.58 2.80 3.58
                 2.80 4.22 4.20 4.22 ;
        RECT  2.96 1.44 3.96 1.76 ;
        POLYGON  1.88 2.08 0.18 2.08 0.18 1.44 0.50 1.44 0.50 1.76 1.56 1.76
                 1.56 1.44 1.88 1.44 ;
    END
END ao22_2

MACRO ao22_1
    CLASS CORE ;
    FOREIGN ao22_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.76 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.45  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.48 2.72 1.12 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.45  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.40 1.76 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.45  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.40 2.72 3.04 3.04 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.45  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.40 4.32 3.04 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  5.60 4.54 5.26 4.54 5.26 4.22 5.28 4.22 5.28 2.09 5.26 2.09
                 5.26 1.77 5.60 1.77 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  5.76 0.90 4.84 0.90 4.84 1.76 4.52 1.76 4.52 0.90 1.20 0.90
                 1.20 1.30 0.88 1.30 0.88 0.90 0.00 0.90 0.00 -0.90 5.76 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.76 6.66 0.00 6.66 0.00 4.86 1.10 4.86 1.10 4.58 1.42 4.58
                 1.42 4.86 4.56 4.86 4.56 4.22 4.88 4.22 4.88 4.86 5.76 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.94 3.90 3.18 3.90 3.18 3.58 3.36 3.58 3.36 2.40 2.26 2.40
                 2.26 1.74 2.58 1.74 2.58 2.08 3.68 2.08 3.68 3.58 4.62 3.58
                 4.62 3.34 4.94 3.34 ;
        POLYGON  4.20 4.54 1.80 4.54 1.80 3.90 0.72 3.90 0.72 4.54 0.40 4.54
                 0.40 3.58 2.12 3.58 2.12 4.22 4.20 4.22 ;
        RECT  2.96 1.44 3.96 1.76 ;
        POLYGON  1.88 2.08 0.18 2.08 0.18 1.44 0.50 1.44 0.50 1.76 1.56 1.76
                 1.56 1.44 1.88 1.44 ;
    END
END ao22_1

MACRO ao222_4
    CLASS CORE ;
    FOREIGN ao222_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.96 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.92 2.58 6.24 3.22 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.58 4.96 3.22 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.58 3.04 3.22 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.58 4.32 3.22 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.58 1.76 3.22 ;
        END
    END e
    PIN f
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.58 0.48 3.22 ;
        END
    END f
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.77  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.80 3.04 8.38 3.04 8.38 4.54 8.06 4.54 8.06 3.90 6.98 3.90
                 6.98 4.54 6.66 4.54 6.66 3.58 8.06 3.58 8.06 1.54 7.12 1.54
                 7.12 1.22 8.38 1.22 8.38 2.72 8.80 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.96 0.90 6.74 0.90 6.74 1.54 6.42 1.54 6.42 0.90 2.58 0.90
                 2.58 1.54 2.26 1.54 2.26 0.90 0.00 0.90 0.00 -0.90 8.96 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  8.96 6.66 0.00 6.66 0.00 4.86 5.28 4.86 5.28 4.22 5.60 4.22
                 5.60 4.86 7.36 4.86 7.36 4.22 7.68 4.22 7.68 4.86 8.96 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  7.35 2.92 7.03 2.92 7.03 2.18 2.40 2.18 2.40 3.86 1.12 3.86
                 1.12 3.54 2.08 3.54 2.08 2.18 0.18 2.18 0.18 1.22 0.50 1.22
                 0.50 1.86 4.34 1.86 4.34 1.22 4.66 1.22 4.66 1.86 7.35 1.86 ;
        POLYGON  6.30 4.54 5.98 4.54 5.98 3.86 4.90 3.86 4.90 4.54 4.58 4.54
                 4.58 3.86 3.20 3.86 3.20 3.54 6.30 3.54 ;
        RECT  5.04 1.22 6.04 1.54 ;
        POLYGON  4.22 4.54 0.42 4.54 0.42 3.54 0.74 3.54 0.74 4.22 4.22 4.22 ;
        RECT  2.96 1.22 3.96 1.54 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END ao222_4

MACRO ao222_2
    CLASS CORE ;
    FOREIGN ao222_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.32 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.92 2.58 6.24 3.22 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.58 4.96 3.22 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.62 3.04 3.26 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.58 4.32 3.22 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.58 1.76 3.22 ;
        END
    END e
    PIN f
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.58 0.48 3.22 ;
        END
    END f
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.16 3.04 8.00 3.04 8.00 4.54 7.68 4.54 7.68 1.54 7.36 1.54
                 7.36 1.22 8.00 1.22 8.00 2.72 8.16 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 0.90 2.58 0.90 2.58 1.54 2.26 1.54 2.26 0.90 0.00 0.90
                 0.00 -0.90 8.32 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 6.66 0.00 6.66 0.00 4.86 5.60 4.86 5.60 4.22 5.92 4.22
                 5.92 4.86 6.98 4.86 6.98 4.22 7.30 4.22 7.30 4.86 8.32 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  7.35 3.04 7.03 3.04 7.03 2.18 2.40 2.18 2.40 3.86 1.20 3.86
                 1.20 3.54 2.08 3.54 2.08 2.18 0.18 2.18 0.18 1.22 0.50 1.22
                 0.50 1.86 4.34 1.86 4.34 1.22 4.66 1.22 4.66 1.86 7.35 1.86 ;
        POLYGON  6.62 4.54 6.30 4.54 6.30 3.86 5.22 3.86 5.22 4.54 4.90 4.54
                 4.90 3.86 3.44 3.86 3.44 3.54 6.62 3.54 ;
        RECT  5.04 1.22 6.04 1.54 ;
        POLYGON  4.54 4.54 0.42 4.54 0.42 3.54 0.74 3.54 0.74 4.22 4.54 4.22 ;
        RECT  2.96 1.22 3.96 1.54 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END ao222_2

MACRO ao222_1
    CLASS CORE ;
    FOREIGN ao222_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.32 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.92 2.72 6.56 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.72 5.28 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.36 3.04 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.68 2.72 4.32 3.04 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.12 2.72 1.76 3.04 ;
        END
    END e
    PIN f
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.72 0.80 3.04 ;
        END
    END f
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.16 3.04 8.00 3.04 8.00 4.54 7.68 4.54 7.68 1.54 7.36 1.54
                 7.36 1.22 8.00 1.22 8.00 2.72 8.16 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 0.90 6.85 0.90 6.85 1.54 6.53 1.54 6.53 0.90 2.58 0.90
                 2.58 1.54 2.26 1.54 2.26 0.90 0.00 0.90 0.00 -0.90 8.32 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 6.66 0.00 6.66 0.00 4.86 6.98 4.86 6.98 4.22 7.30 4.22
                 7.30 4.86 8.32 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  7.35 3.04 7.03 3.04 7.03 2.18 2.40 2.18 2.40 3.86 1.20 3.86
                 1.20 3.54 2.08 3.54 2.08 2.18 0.18 2.18 0.18 1.22 0.50 1.22
                 0.50 1.86 4.34 1.86 4.34 1.22 4.66 1.22 4.66 1.86 7.35 1.86 ;
        POLYGON  6.62 4.54 4.90 4.54 4.90 3.86 3.44 3.86 3.44 3.54 5.22 3.54
                 5.22 4.22 6.62 4.22 ;
        RECT  5.04 1.22 6.04 1.54 ;
        RECT  0.42 4.22 4.54 4.54 ;
        RECT  2.96 1.22 3.96 1.54 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END ao222_1

MACRO ao221_4
    CLASS CORE ;
    FOREIGN ao221_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  7.02 2.62 7.52 3.06 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.92 2.08 6.56 2.44 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  2.76 2.58 2.44 2.58 2.44 2.40 2.08 2.40 2.08 2.08 2.76 2.08 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.24 3.36 5.88 3.68 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.39 2.62 1.76 3.18 ;
        END
    END e
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  0.52 1.54 0.48 1.54 0.48 4.22 0.52 4.22 0.52 4.54 0.16 4.54
                 0.16 1.22 0.52 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 7.68 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 6.66 0.00 6.66 0.00 4.86 0.90 4.86 0.90 4.22 1.22 4.22
                 1.22 4.86 7.68 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  5.76 1.22 7.46 1.54 ;
        POLYGON  7.46 4.54 2.28 4.54 2.28 4.22 7.14 4.22 7.14 3.58 7.46 3.58 ;
        POLYGON  5.38 1.54 5.32 1.54 5.32 2.46 4.92 2.86 4.92 3.86 2.96 3.86
                 2.96 3.54 4.60 3.54 4.60 2.72 5.00 2.32 5.00 1.54 1.44 1.54
                 1.44 2.12 1.12 2.12 1.12 2.44 0.80 2.44 0.80 1.80 1.12 1.80
                 1.12 1.22 5.38 1.22 ;
        RECT  3.08 1.86 4.68 2.18 ;
        POLYGON  3.98 3.22 2.64 3.22 2.64 3.86 1.90 3.86 1.90 4.54 1.58 4.54
                 1.58 3.54 2.32 3.54 2.32 2.90 3.98 2.90 ;
    END
END ao221_4

MACRO ao221_2
    CLASS CORE ;
    FOREIGN ao221_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  7.02 2.62 7.52 3.06 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.92 2.08 6.56 2.44 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  2.76 2.58 2.08 2.58 2.08 2.08 2.40 2.08 2.40 2.26 2.76 2.26 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.24 3.36 5.88 3.68 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.50 1.76 3.14 ;
        END
    END e
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  0.52 1.54 0.48 1.54 0.48 4.22 0.52 4.22 0.52 4.54 0.16 4.54
                 0.16 1.22 0.52 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 7.68 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 6.66 0.00 6.66 0.00 4.86 0.90 4.86 0.90 4.22 1.22 4.22
                 1.22 4.86 7.68 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  5.76 1.22 7.46 1.54 ;
        POLYGON  7.46 4.54 2.28 4.54 2.28 4.22 7.14 4.22 7.14 3.58 7.46 3.58 ;
        POLYGON  5.38 1.54 5.32 1.54 5.32 2.46 4.88 2.90 4.88 3.54 4.92 3.54
                 4.92 3.86 2.96 3.86 2.96 3.54 4.56 3.54 4.56 2.76 5.00 2.32
                 5.00 1.54 1.44 1.54 1.44 2.02 0.80 2.02 0.80 1.70 1.12 1.70
                 1.12 1.22 5.38 1.22 ;
        RECT  3.08 1.86 4.68 2.18 ;
        POLYGON  3.98 3.22 2.64 3.22 2.64 3.86 1.90 3.86 1.90 4.54 1.58 4.54
                 1.58 3.54 2.32 3.54 2.32 2.90 3.98 2.90 ;
    END
END ao221_2

MACRO ao221_1
    CLASS CORE ;
    FOREIGN ao221_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.04 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.62 1.12 3.36 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.66 0.48 3.40 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.50 1.92 3.04 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.50  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.50 4.96 3.24 ;
        END
    END d
    PIN e
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 2.72 5.71 3.24 ;
        END
    END e
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  6.88 3.68 6.74 3.68 6.74 4.54 6.42 4.54 6.42 1.22 6.74 1.22
                 6.74 3.36 6.88 3.36 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  7.04 0.90 6.04 0.90 6.04 1.54 5.04 1.54 5.04 0.90 2.58 0.90
                 2.58 1.54 2.26 1.54 2.26 0.90 0.00 0.90 0.00 -0.90 7.04 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.04 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.50 1.20 4.50
                 1.20 4.86 5.72 4.86 5.72 4.44 6.04 4.44 6.04 4.86 7.04 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  6.06 2.40 5.74 2.40 5.74 2.18 3.68 2.18 3.68 2.92 3.98 2.92
                 3.98 3.24 2.26 3.24 2.26 2.92 3.36 2.92 3.36 2.18 0.18 2.18
                 0.18 1.22 0.50 1.22 0.50 1.86 4.34 1.86 4.34 1.22 4.66 1.22
                 4.66 1.86 6.06 1.86 ;
        POLYGON  5.36 4.54 5.04 4.54 5.04 3.88 1.90 3.88 1.90 4.18 0.50 4.18
                 0.50 4.54 0.18 4.54 0.18 3.86 1.58 3.86 1.58 3.56 5.36 3.56 ;
        RECT  2.96 4.22 4.66 4.54 ;
        RECT  2.96 1.22 3.96 1.54 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END ao221_1

MACRO ao21_4
    CLASS CORE ;
    FOREIGN ao21_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.48 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.08 4.32 2.72 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.08 3.04 2.72 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.72 1.86 3.26 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  0.52 1.54 0.48 1.54 0.48 4.22 0.52 4.22 0.52 4.54 0.16 4.54
                 0.16 1.22 0.52 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  4.48 0.90 3.54 0.90 3.54 1.12 3.22 1.12 3.22 0.90 0.00 0.90
                 0.00 -0.90 4.48 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  4.48 6.66 0.00 6.66 0.00 4.86 1.02 4.86 1.02 4.22 1.34 4.22
                 1.34 4.86 4.48 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.24 1.76 2.54 1.76 2.54 1.22 2.86 1.22 2.86 1.44 3.92 1.44
                 3.92 1.22 4.24 1.22 ;
        POLYGON  4.24 4.32 3.92 4.32 3.92 3.90 0.80 3.90 0.80 1.98 1.84 1.98
                 1.84 1.22 2.16 1.22 2.16 2.30 1.12 2.30 1.12 3.58 4.24 3.58 ;
        RECT  1.84 4.22 3.54 4.54 ;
    END
END ao21_4

MACRO ao21_2
    CLASS CORE ;
    FOREIGN ao21_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.48 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.08 4.32 2.72 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.14 3.04 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.62 1.76 3.26 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  0.52 1.54 0.48 1.54 0.48 4.22 0.52 4.22 0.52 4.54 0.16 4.54
                 0.16 1.22 0.52 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  4.48 0.90 3.44 0.90 3.44 1.12 3.12 1.12 3.12 0.90 1.28 0.90
                 1.28 1.54 0.96 1.54 0.96 0.90 0.00 0.90 0.00 -0.90 4.48 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 4.48 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.14 1.76 2.44 1.76 2.44 1.22 2.76 1.22 2.76 1.44 3.82 1.44
                 3.82 1.22 4.14 1.22 ;
        POLYGON  4.14 4.32 3.82 4.32 3.82 3.90 0.80 3.90 0.80 1.98 1.74 1.98
                 1.74 1.22 2.06 1.22 2.06 2.30 1.12 2.30 1.12 3.58 4.14 3.58 ;
        RECT  1.74 4.22 3.44 4.54 ;
    END
END ao21_2

MACRO ao21_1
    CLASS CORE ;
    FOREIGN ao21_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.48 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.08 4.32 2.72 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.08 3.04 2.72 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.72 1.86 3.26 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  0.52 1.54 0.48 1.54 0.48 4.22 0.52 4.22 0.52 4.54 0.16 4.54
                 0.16 1.22 0.52 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  4.48 0.90 3.54 0.90 3.54 1.12 3.22 1.12 3.22 0.90 1.31 0.90
                 1.31 1.54 0.99 1.54 0.99 0.90 0.00 0.90 0.00 -0.90 4.48 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  4.48 6.66 0.00 6.66 0.00 4.86 0.99 4.86 0.99 4.28 1.31 4.28
                 1.31 4.86 4.48 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.24 1.76 2.54 1.76 2.54 1.22 2.86 1.22 2.86 1.44 3.92 1.44
                 3.92 1.22 4.24 1.22 ;
        POLYGON  4.24 4.32 3.92 4.32 3.92 3.90 0.80 3.90 0.80 1.98 1.84 1.98
                 1.84 1.22 2.16 1.22 2.16 2.30 1.12 2.30 1.12 3.58 4.24 3.58 ;
        RECT  1.84 4.22 3.54 4.54 ;
    END
END ao21_1

MACRO ao211_4
    CLASS CORE ;
    FOREIGN ao211_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.76 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.50 1.76 3.24 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.50 0.48 3.24 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.50 4.32 3.24 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.50 3.04 3.24 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  5.60 4.54 5.26 4.54 5.26 4.22 5.28 4.22 5.28 1.54 5.26 1.54
                 5.26 1.22 5.60 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  5.76 0.90 4.66 0.90 4.66 1.54 4.34 1.54 4.34 0.90 2.58 0.90
                 2.58 1.54 2.26 1.54 2.26 0.90 0.00 0.90 0.00 -0.90 5.76 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.76 6.66 0.00 6.66 0.00 4.86 4.44 4.86 4.44 3.58 4.76 3.58
                 4.76 4.86 5.76 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.96 2.44 4.64 2.44 4.64 2.18 1.12 2.18 1.12 3.58 1.90 3.58
                 1.90 3.90 0.50 3.90 0.50 4.54 0.18 4.54 0.18 3.58 0.80 3.58
                 0.80 2.18 0.18 2.18 0.18 1.22 0.50 1.22 0.50 1.86 2.96 1.86
                 2.96 1.22 3.84 1.22 3.84 1.86 4.96 1.86 ;
        RECT  2.96 3.58 3.96 4.54 ;
        POLYGON  2.58 4.54 0.88 4.54 0.88 4.22 2.26 4.22 2.26 3.58 2.58 3.58 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END ao211_4

MACRO ao211_2
    CLASS CORE ;
    FOREIGN ao211_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.50 1.76 3.24 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.50 0.48 3.24 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.50 4.32 3.24 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.50 3.04 3.24 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 1.22 5.60 4.54 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 0.90 4.66 0.90 4.66 1.54 4.34 1.54 4.34 0.90 2.58 0.90
                 2.58 1.54 2.26 1.54 2.26 0.90 0.00 0.90 0.00 -0.90 6.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 6.66 0.00 6.66 0.00 4.86 4.47 4.86 4.47 4.22 4.79 4.22
                 4.79 4.86 6.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.96 2.44 4.64 2.44 4.64 2.18 1.12 2.18 1.12 3.58 1.90 3.58
                 1.90 3.90 0.50 3.90 0.50 4.54 0.18 4.54 0.18 3.58 0.80 3.58
                 0.80 2.18 0.18 2.18 0.18 1.22 0.50 1.22 0.50 1.86 2.96 1.86
                 2.96 1.22 3.84 1.22 3.84 1.86 4.96 1.86 ;
        RECT  2.96 3.58 3.96 4.54 ;
        POLYGON  2.58 4.54 0.88 4.54 0.88 4.22 2.26 4.22 2.26 3.58 2.58 3.58 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END ao211_2

MACRO ao211_1
    CLASS CORE ;
    FOREIGN ao211_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.50 1.76 3.24 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.16 2.50 0.48 3.24 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.00 2.50 4.32 3.24 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.50 3.04 3.24 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.28 1.22 5.60 4.54 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 0.90 4.66 0.90 4.66 1.54 4.34 1.54 4.34 0.90 2.58 0.90
                 2.58 1.54 2.26 1.54 2.26 0.90 0.00 0.90 0.00 -0.90 6.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 6.66 0.00 6.66 0.00 4.86 4.46 4.86 4.46 4.22 4.78 4.22
                 4.78 4.86 6.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.96 2.44 4.64 2.44 4.64 2.18 1.12 2.18 1.12 3.58 1.90 3.58
                 1.90 3.90 0.50 3.90 0.50 4.54 0.18 4.54 0.18 3.58 0.80 3.58
                 0.80 2.18 0.18 2.18 0.18 1.22 0.50 1.22 0.50 1.86 2.96 1.86
                 2.96 1.22 3.86 1.22 3.86 1.86 4.96 1.86 ;
        POLYGON  3.96 4.54 2.96 4.54 2.96 4.22 3.64 4.22 3.64 3.58 3.96 3.58 ;
        RECT  0.88 4.22 2.58 4.54 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END ao211_1

MACRO and4_8
    CLASS CORE ;
    FOREIGN and4_8 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.08 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.22  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.60 1.12 3.24 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.04 3.39 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.22  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  5.08 2.64 5.72 3.04 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.15  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.72 4.26 3.16 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.46  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  13.86 1.54 12.96 1.54 12.96 2.08 13.28 2.08 13.28 2.40
                 12.96 2.40 12.96 3.90 12.64 3.90 12.64 3.26 11.56 3.26
                 11.56 3.90 11.24 3.90 11.24 2.94 12.64 2.94 12.64 1.54
                 7.94 1.54 7.94 1.22 13.86 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  14.08 0.90 4.04 0.90 4.04 1.54 3.72 1.54 3.72 0.90 0.00 0.90
                 0.00 -0.90 14.08 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  14.08 6.66 0.00 6.66 0.00 4.86 8.46 4.86 8.46 4.22 8.78 4.22
                 8.78 4.86 14.08 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  13.66 4.54 9.16 4.54 9.16 3.90 8.02 3.90 8.02 4.54 7.70 4.54
                 7.70 3.58 9.48 3.58 9.48 4.22 10.54 4.22 10.54 3.58 10.86 3.58
                 10.86 4.22 11.94 4.22 11.94 3.58 12.26 3.58 12.26 4.22
                 13.34 4.22 13.34 3.58 13.66 3.58 ;
        POLYGON  11.98 2.58 9.52 2.58 9.52 3.26 7.38 3.26 7.38 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.86 1.90 1.86 1.90 2.18 0.48 2.18
                 0.48 4.22 7.06 4.22 7.06 2.94 9.20 2.94 9.20 2.26 11.98 2.26 ;
        POLYGON  8.58 2.60 7.26 2.60 7.26 2.18 6.44 2.18 6.44 3.90 4.66 3.90
                 4.66 3.58 6.12 3.58 6.12 2.18 5.80 2.18 5.80 1.86 7.26 1.86
                 7.26 1.22 7.58 1.22 7.58 2.28 8.58 2.28 ;
        RECT  4.42 1.22 6.82 1.54 ;
        RECT  0.88 1.22 3.34 1.54 ;
    END
END and4_8

MACRO and4_4
    CLASS CORE ;
    FOREIGN and4_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.24 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.62 1.76 3.26 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.62 2.40 3.26 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.08 3.88 2.59 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.36 3.04 3.14 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.68  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.64 1.54 8.80 1.54 8.80 2.94 8.94 2.94 8.94 3.90 8.62 3.90
                 8.62 3.26 7.54 3.26 7.54 3.90 7.22 3.90 7.22 2.94 8.48 2.94
                 8.48 1.54 5.06 1.54 5.06 1.22 9.64 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  10.24 0.90 2.58 0.90 2.58 1.54 2.26 1.54 2.26 0.90 0.00 0.90
                 0.00 -0.90 10.24 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 10.24 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  9.64 4.54 5.13 4.54 5.13 4.22 7.92 4.22 7.92 3.58 8.24 3.58
                 8.24 4.22 9.32 4.22 9.32 3.58 9.64 3.58 ;
        POLYGON  7.96 2.59 6.12 2.59 6.12 3.90 4.81 3.90 4.81 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.56 0.48 1.56 0.48 4.22 4.49 4.22
                 4.49 3.58 5.80 3.58 5.80 2.27 7.96 2.27 ;
        POLYGON  5.12 2.53 4.66 2.53 4.66 3.26 4.16 3.26 4.16 3.90 3.44 3.90
                 3.44 3.58 3.84 3.58 3.84 2.94 4.34 2.94 4.34 1.22 4.66 1.22
                 4.66 2.21 5.12 2.21 ;
        RECT  2.96 1.22 3.96 1.54 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END and4_4

MACRO and4_2
    CLASS CORE ;
    FOREIGN and4_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.32 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.60 1.12 3.24 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.72 1.76 3.39 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.58  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.44 2.46 3.04 2.46 3.04 2.40 2.72 2.40 2.72 2.08 3.44 2.08 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.58  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.72 2.74 3.16 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.85  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.16 3.26 7.94 3.26 7.94 4.54 7.62 4.54 7.62 3.26 6.54 3.26
                 6.54 3.90 6.22 3.90 6.22 2.94 7.84 2.94 7.84 1.56 5.02 1.56
                 5.02 1.24 8.16 1.24 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 0.90 2.58 0.90 2.58 1.54 2.26 1.54 2.26 0.90 0.00 0.90
                 0.00 -0.90 8.32 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 8.32 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  7.24 4.54 4.84 4.54 4.84 4.22 6.92 4.22 6.92 3.58 7.24 3.58 ;
        POLYGON  6.96 2.62 5.46 2.62 5.46 3.90 4.52 3.90 4.52 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.56 0.48 1.56 0.48 4.22 4.20 4.22
                 4.20 3.58 5.14 3.58 5.14 2.30 6.96 2.30 ;
        POLYGON  4.82 2.60 4.08 2.60 4.08 3.10 3.52 3.10 3.52 3.90 3.20 3.90
                 3.20 2.78 3.76 2.78 3.76 2.28 4.34 2.28 4.34 1.22 4.66 1.22
                 4.66 2.28 4.82 2.28 ;
        RECT  2.96 1.22 3.96 1.54 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END and4_2

MACRO and4_1
    CLASS CORE ;
    FOREIGN and4_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.04 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.60 1.12 3.24 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.72 1.76 3.39 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.58  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.44 2.46 3.04 2.46 3.04 2.40 2.72 2.40 2.72 2.08 3.44 2.08 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.58  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.72 2.74 3.16 ;
        END
    END d
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.13  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  6.74 1.54 6.54 1.54 6.54 4.54 6.22 4.54 6.22 2.40 5.92 2.40
                 5.92 2.08 6.22 2.08 6.22 1.54 5.02 1.54 5.02 1.22 6.74 1.22 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  7.04 0.90 2.58 0.90 2.58 1.54 2.26 1.54 2.26 0.90 0.00 0.90
                 0.00 -0.90 7.04 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
        RECT  0.00 4.86 7.04 6.66 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  4.84 4.22 5.84 4.54 ;
        POLYGON  5.56 2.62 5.46 2.62 5.46 3.90 4.52 3.90 4.52 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.56 0.48 1.56 0.48 4.22 4.20 4.22
                 4.20 3.58 5.14 3.58 5.14 2.30 5.56 2.30 ;
        POLYGON  4.82 2.60 4.08 2.60 4.08 3.10 3.52 3.10 3.52 3.90 3.20 3.90
                 3.20 2.78 3.76 2.78 3.76 2.28 4.34 2.28 4.34 1.22 4.66 1.22
                 4.66 2.28 4.82 2.28 ;
        RECT  2.96 1.22 3.96 1.54 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END and4_1

MACRO and3_8
    CLASS CORE ;
    FOREIGN and3_8 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 10.24 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.98  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.18 2.72 1.76 3.37 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.98  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.12 3.37 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.98  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  4.64 2.72 5.04 3.37 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.29  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  9.62 1.96 8.22 1.96 8.22 3.78 9.30 3.78 9.30 3.10 9.62 3.10
                 9.62 4.10 6.50 4.10 6.50 3.16 6.82 3.16 6.82 3.78 7.90 3.78
                 7.90 3.04 7.84 3.04 7.84 2.72 7.90 2.72 7.90 1.96 6.50 1.96
                 6.50 1.64 9.62 1.64 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  10.24 0.90 8.92 0.90 8.92 1.32 8.60 1.32 8.60 0.90 7.52 0.90
                 7.52 1.32 7.20 1.32 7.20 0.90 0.00 0.90 0.00 -0.90 10.24 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  10.24 6.66 0.00 6.66 0.00 4.86 7.20 4.86 7.20 4.42 7.52 4.42
                 7.52 4.86 8.60 4.86 8.60 4.42 8.92 4.42 8.92 4.86 10.24 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  7.44 2.66 6.14 2.66 6.14 4.54 0.18 4.54 0.18 1.22 0.50 1.22
                 0.50 1.86 1.98 1.86 1.98 2.18 0.50 2.18 0.50 4.22 5.82 4.22
                 5.82 2.34 7.44 2.34 ;
        RECT  3.04 1.22 6.14 1.54 ;
        POLYGON  4.14 2.18 2.34 2.18 2.34 1.54 0.88 1.54 0.88 1.22 2.66 1.22
                 2.66 1.86 4.14 1.86 ;
    END
END and3_8

MACRO and3_4
    CLASS CORE ;
    FOREIGN and3_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 3.26 1.50 3.68 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.40 2.40 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.08 3.36 2.43 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.97  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.96 3.04 4.90 3.04 4.90 4.54 4.58 4.54 4.58 1.30 4.90 1.30
                 4.90 2.72 4.96 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 0.90 5.60 0.90 5.60 1.08 5.28 1.08 5.28 0.90 4.06 0.90
                 4.06 1.08 3.74 1.08 3.74 0.90 0.00 0.90 0.00 -0.90 6.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 6.66 0.00 6.66 0.00 4.86 1.20 4.86 1.20 4.68 1.52 4.68
                 1.52 4.86 3.75 4.86 3.75 4.28 4.07 4.28 4.07 4.86 5.28 4.86
                 5.28 4.28 5.60 4.28 5.60 4.86 6.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.12 3.09 3.26 3.09 3.26 4.36 0.16 4.36 0.16 1.22 0.50 1.22
                 0.50 1.54 0.48 1.54 0.48 4.04 2.94 4.04 2.94 2.77 3.80 2.77
                 3.80 2.59 4.12 2.59 ;
        RECT  2.26 1.22 3.26 1.54 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END and3_4

MACRO and3_2
    CLASS CORE ;
    FOREIGN and3_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 3.26 1.50 3.68 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.40 2.40 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.08 3.36 2.43 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.96 3.04 4.90 3.04 4.90 4.54 4.58 4.54 4.58 1.30 4.90 1.30
                 4.90 2.72 4.96 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 0.90 4.06 0.90 4.06 1.08 3.74 1.08 3.74 0.90 0.00 0.90
                 0.00 -0.90 5.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 6.66 0.00 6.66 0.00 4.86 1.20 4.86 1.20 4.68 1.52 4.68
                 1.52 4.86 3.75 4.86 3.75 4.28 4.07 4.28 4.07 4.86 5.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.12 3.09 3.26 3.09 3.26 4.36 0.16 4.36 0.16 1.22 0.50 1.22
                 0.50 1.54 0.48 1.54 0.48 4.04 2.94 4.04 2.94 2.77 3.80 2.77
                 3.80 2.59 4.12 2.59 ;
        RECT  2.26 1.22 3.26 1.54 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END and3_2

MACRO and3_1
    CLASS CORE ;
    FOREIGN and3_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 3.26 1.50 3.68 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.40 2.40 3.04 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.49  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.72 2.72 3.36 3.04 ;
        END
    END c
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.96 3.04 4.90 3.04 4.90 4.54 4.58 4.54 4.58 1.22 4.90 1.22
                 4.90 2.72 4.96 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 0.90 4.06 0.90 4.06 1.08 3.74 1.08 3.74 0.90 0.00 0.90
                 0.00 -0.90 5.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 6.66 0.00 6.66 0.00 4.86 1.20 4.86 1.20 4.68 1.52 4.68
                 1.52 4.86 3.75 4.86 3.75 4.28 4.07 4.28 4.07 4.86 5.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.12 3.68 3.26 3.68 3.26 4.36 0.16 4.36 0.16 1.22 0.50 1.22
                 0.50 1.54 0.48 1.54 0.48 4.04 2.94 4.04 2.94 3.36 3.80 3.36
                 3.80 3.26 4.12 3.26 ;
        RECT  2.26 1.22 3.26 1.54 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END and3_1

MACRO and2a_8
    CLASS CORE ;
    FOREIGN and2a_8 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.60 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.45  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.72 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.13  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.78 2.72 4.42 3.04 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.29  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  8.86 1.96 7.46 1.96 7.46 2.72 7.52 2.72 7.52 3.04 7.46 3.04
                 7.46 3.78 8.54 3.78 8.54 3.10 8.86 3.10 8.86 4.10 5.74 4.10
                 5.74 3.16 6.06 3.16 6.06 3.78 7.14 3.78 7.14 1.96 5.74 1.96
                 5.74 1.64 8.86 1.64 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  9.60 0.90 8.16 0.90 8.16 1.32 7.84 1.32 7.84 0.90 6.76 0.90
                 6.76 1.32 6.44 1.32 6.44 0.90 4.67 0.90 4.67 1.08 4.35 1.08
                 4.35 0.90 1.20 0.90 1.20 1.66 0.88 1.66 0.88 0.90 0.00 0.90
                 0.00 -0.90 9.60 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  9.60 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.66 1.20 4.66
                 1.20 4.86 2.26 4.86 2.26 4.68 2.58 4.68 2.58 4.86 4.35 4.86
                 4.35 4.68 4.67 4.68 4.67 4.86 6.44 4.86 6.44 4.42 6.76 4.42
                 6.76 4.86 7.84 4.86 7.84 4.42 8.16 4.42 8.16 4.86 9.60 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  6.68 2.66 5.38 2.66 5.38 4.37 5.06 4.37 5.06 4.36 1.54 4.36
                 1.54 4.04 2.18 4.04 2.18 2.83 1.54 2.83 1.54 1.22 3.28 1.22
                 3.28 1.54 1.86 1.54 1.86 2.51 2.50 2.51 2.50 4.04 5.06 4.04
                 5.06 2.34 6.68 2.34 ;
        POLYGON  5.38 1.72 3.92 1.72 3.92 2.18 2.26 2.18 2.26 1.86 3.60 1.86
                 3.60 1.40 5.38 1.40 ;
        POLYGON  1.78 3.58 0.48 3.58 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 3.26 1.78 3.26 ;
    END
END and2a_8

MACRO and2a_4
    CLASS CORE ;
    FOREIGN and2a_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 6.40 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.45  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.72 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.03 3.22 3.68 3.68 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.97  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.96 3.04 4.90 3.04 4.90 4.54 4.58 4.54 4.58 1.64 4.90 1.64
                 4.90 2.72 4.96 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 0.90 5.60 0.90 5.60 1.08 5.28 1.08 5.28 0.90 4.06 0.90
                 4.06 1.08 3.74 1.08 3.74 0.90 0.00 0.90 0.00 -0.90 6.40 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  6.40 6.66 0.00 6.66 0.00 4.86 3.75 4.86 3.75 4.22 4.07 4.22
                 4.07 4.86 5.28 4.86 5.28 4.22 5.60 4.22 5.60 4.86 6.40 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.12 2.90 2.58 2.90 2.58 4.22 3.26 4.22 3.26 4.54 1.56 4.54
                 1.56 4.22 2.26 4.22 2.26 2.18 1.56 2.18 1.56 1.22 1.88 1.22
                 1.88 1.86 2.58 1.86 2.58 2.58 4.12 2.58 ;
        RECT  2.26 1.22 3.26 1.54 ;
        POLYGON  1.36 3.58 0.48 3.58 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 3.26 1.36 3.26 ;
    END
END and2a_4

MACRO and2a_2
    CLASS CORE ;
    FOREIGN and2a_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.45  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.72 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.03 3.22 3.68 3.68 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.96 3.04 4.90 3.04 4.90 4.54 4.58 4.54 4.58 1.64 4.90 1.64
                 4.90 2.72 4.96 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 0.90 4.06 0.90 4.06 1.08 3.74 1.08 3.74 0.90 0.00 0.90
                 0.00 -0.90 5.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 6.66 0.00 6.66 0.00 4.86 3.75 4.86 3.75 4.22 4.07 4.22
                 4.07 4.86 5.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.12 2.90 2.58 2.90 2.58 4.22 3.26 4.22 3.26 4.54 1.56 4.54
                 1.56 4.22 2.26 4.22 2.26 2.18 1.56 2.18 1.56 1.22 1.88 1.22
                 1.88 1.86 2.58 1.86 2.58 2.58 4.12 2.58 ;
        RECT  2.26 1.22 3.26 1.54 ;
        POLYGON  1.36 3.58 0.48 3.58 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 3.26 1.36 3.26 ;
    END
END and2a_2

MACRO and2a_1
    CLASS CORE ;
    FOREIGN and2a_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.45  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.08 1.12 2.72 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.04 3.68 2.68 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.96 3.04 4.90 3.04 4.90 4.37 4.58 4.37 4.58 1.22 4.90 1.22
                 4.90 2.72 4.96 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 0.90 4.06 0.90 4.06 1.08 3.74 1.08 3.74 0.90 0.00 0.90
                 0.00 -0.90 5.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 6.66 0.00 6.66 0.00 4.86 3.75 4.86 3.75 4.68 4.07 4.68
                 4.07 4.86 5.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  4.12 3.68 3.54 3.68 3.54 4.36 1.54 4.36 1.54 4.04 2.26 4.04
                 2.26 2.18 1.56 2.18 1.56 1.22 1.88 1.22 1.88 1.86 2.58 1.86
                 2.58 4.04 3.22 4.04 3.22 3.36 3.80 3.36 3.80 3.26 4.12 3.26 ;
        RECT  2.26 1.22 3.26 1.54 ;
        POLYGON  1.36 3.58 0.48 3.58 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.22 0.50 1.22 0.50 1.54 0.48 1.54 0.48 3.26 1.36 3.26 ;
    END
END and2a_1

MACRO and2_8
    CLASS CORE ;
    FOREIGN and2_8 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.32 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.13  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.06 3.26 1.76 3.68 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.13  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 3.00 3.68 3.68 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.31  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.72 3.68 4.60 3.68 4.60 3.36 7.40 3.36 7.40 1.95 4.60 1.95
                 4.60 1.63 7.72 1.63 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 0.90 7.02 0.90 7.02 1.30 6.70 1.30 6.70 0.90 5.62 0.90
                 5.62 1.31 5.30 1.31 5.30 0.90 0.00 0.90 0.00 -0.90 8.32 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  8.32 6.66 0.00 6.66 0.00 4.86 1.12 4.86 1.12 4.68 1.44 4.68
                 1.44 4.86 3.21 4.86 3.21 4.68 3.56 4.68 3.56 4.86 5.30 4.86
                 5.30 4.11 5.63 4.11 5.63 4.86 6.70 4.86 6.70 4.11 7.03 4.11
                 7.03 4.86 8.32 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  6.30 2.68 3.82 2.68 3.82 2.18 0.74 2.18 0.74 4.04 4.24 4.04
                 4.24 4.36 0.42 4.36 0.42 1.86 4.14 1.86 4.14 2.36 6.30 2.36 ;
        RECT  1.12 1.22 4.25 1.54 ;
    END
END and2_8

MACRO and2_4
    CLASS CORE ;
    FOREIGN and2_4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.12 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 2.62 1.12 3.26 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.44 2.62 1.76 3.26 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.33  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.96 3.58 4.66 3.58 4.66 4.14 4.34 4.14 4.34 3.86 3.26 3.86
                 3.26 4.14 2.94 4.14 2.94 3.26 3.26 3.26 3.26 3.54 4.34 3.54
                 4.34 3.26 4.64 3.26 4.64 1.96 2.94 1.96 2.94 1.64 4.96 1.64 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 0.90 3.96 0.90 3.96 1.32 3.64 1.32 3.64 0.90 2.58 0.90
                 2.58 1.54 2.26 1.54 2.26 0.90 0.00 0.90 0.00 -0.90 5.12 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  5.12 6.66 0.00 6.66 0.00 4.86 0.42 4.86 0.42 4.22 0.74 4.22
                 0.74 4.86 1.82 4.86 1.82 4.22 2.14 4.22 2.14 4.86 3.64 4.86
                 3.64 4.42 3.96 4.42 3.96 4.86 5.12 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  3.88 2.66 2.59 2.66 2.59 3.90 1.44 3.90 1.44 4.54 1.12 4.54
                 1.12 3.90 0.16 3.90 0.16 1.22 0.50 1.22 0.50 1.56 0.48 1.56
                 0.48 3.58 2.27 3.58 2.27 2.34 3.88 2.34 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END and2_4

MACRO and2_2
    CLASS CORE ;
    FOREIGN and2_2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.84 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 3.26 1.44 3.68 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  2.13 2.68 1.44 2.68 1.44 2.04 1.78 2.04 1.78 2.36 2.13 2.36 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.68 3.04 3.52 3.04 3.52 4.30 3.20 4.30 3.20 1.64 3.52 1.64
                 3.52 2.72 3.68 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  3.84 0.90 2.68 0.90 2.68 1.08 2.36 1.08 2.36 0.90 0.00 0.90
                 0.00 -0.90 3.84 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  3.84 6.66 0.00 6.66 0.00 4.86 2.37 4.86 2.37 4.68 2.69 4.68
                 2.69 4.86 3.84 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  2.88 4.36 0.16 4.36 0.16 1.22 0.50 1.22 0.50 2.10 0.48 2.10
                 0.48 4.04 2.56 4.04 2.56 2.62 2.88 2.62 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END and2_2

MACRO and2_1
    CLASS CORE ;
    FOREIGN and2_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 3.84 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  0.80 3.26 1.44 3.68 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.57  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  2.08 2.04 2.40 2.68 ;
        END
    END b
    PIN x
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.68 3.04 3.52 3.04 3.52 4.06 3.20 4.06 3.20 1.22 3.52 1.22
                 3.52 2.72 3.68 2.72 ;
        END
    END x
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  3.84 0.90 2.68 0.90 2.68 1.08 2.36 1.08 2.36 0.90 0.00 0.90
                 0.00 -0.90 3.84 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  3.84 6.66 0.00 6.66 0.00 4.86 2.37 4.86 2.37 4.68 2.69 4.68
                 2.69 4.86 3.84 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  2.74 3.68 2.16 3.68 2.16 4.36 0.16 4.36 0.16 1.22 0.50 1.22
                 0.50 2.10 0.48 2.10 0.48 4.04 1.84 4.04 1.84 3.36 2.42 3.36
                 2.42 3.26 2.74 3.26 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END and2_1

MACRO adhalf_1
    CLASS CORE ;
    FOREIGN adhalf_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.84 2.18 1.12 2.18 1.12 2.40 0.80 2.40 0.80 1.86 3.84 1.86 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.94 2.58 2.40 3.04 ;
        END
    END b
    PIN co
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  6.24 2.40 6.02 2.40 6.02 3.42 5.70 3.42 5.70 1.22 6.04 1.22
                 6.04 1.54 6.02 1.54 6.02 2.08 6.24 2.08 ;
        END
    END co
    PIN s
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.89  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.52 4.53 7.18 4.53 7.18 4.21 7.20 4.21 7.20 1.54 7.18 1.54
                 7.18 1.22 7.52 1.22 ;
        END
    END s
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 0.90 6.74 0.90 6.74 1.54 6.42 1.54 6.42 0.90 0.00 0.90
                 0.00 -0.90 7.68 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 6.40 4.86 6.40 4.38 6.72 4.38 6.72 4.86 7.68 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  6.88 4.06 5.30 4.06 5.14 3.90 3.98 3.90 3.98 3.58 5.04 3.58
                 5.04 1.22 5.36 1.22 5.36 3.66 5.44 3.74 6.56 3.74 6.56 2.62
                 6.88 2.62 ;
        RECT  2.26 4.22 5.00 4.54 ;
        POLYGON  4.66 1.66 4.34 1.66 4.34 1.54 2.96 1.54 2.96 1.22 4.66 1.22 ;
        POLYGON  3.44 2.92 3.04 2.92 3.04 3.90 1.90 3.90 1.90 4.54 1.58 4.54
                 1.58 3.90 0.48 3.90 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.32 0.50 1.32 0.50 1.64 0.48 1.64 0.48 3.58 2.72 3.58
                 2.72 2.60 3.44 2.60 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END adhalf_1

MACRO adhalf_0
    CLASS CORE ;
    FOREIGN adhalf_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.68 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  3.84 2.18 1.12 2.18 1.12 2.40 0.80 2.40 0.80 1.86 3.84 1.86 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.09  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  1.94 2.58 2.40 3.04 ;
        END
    END b
    PIN co
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.56  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  6.24 2.40 6.02 2.40 6.02 3.42 5.62 3.42 5.62 3.10 5.70 3.10
                 5.70 1.22 6.04 1.22 6.04 1.54 6.02 1.54 6.02 2.08 6.24 2.08 ;
        END
    END co
    PIN s
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.36  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  7.52 4.53 7.18 4.53 7.18 4.21 7.20 4.21 7.20 1.54 7.18 1.54
                 7.18 1.22 7.52 1.22 ;
        END
    END s
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
        RECT  0.00 -0.90 7.68 0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  7.68 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 6.40 4.86 6.40 4.38 6.72 4.38 6.72 4.86 7.68 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  6.88 4.06 5.30 4.06 5.14 3.90 3.98 3.90 3.98 3.58 4.96 3.58
                 4.96 1.98 5.04 1.98 5.04 1.22 5.36 1.22 5.36 2.30 5.28 2.30
                 5.28 3.58 5.44 3.74 6.56 3.74 6.56 2.62 6.88 2.62 ;
        RECT  2.26 4.22 5.00 4.54 ;
        POLYGON  4.66 1.66 4.34 1.66 4.34 1.54 2.96 1.54 2.96 1.22 4.66 1.22 ;
        POLYGON  3.44 2.92 3.04 2.92 3.04 3.90 1.90 3.90 1.90 4.54 1.58 4.54
                 1.58 3.90 0.48 3.90 0.48 4.22 0.50 4.22 0.50 4.54 0.16 4.54
                 0.16 1.32 0.50 1.32 0.50 1.64 0.48 1.64 0.48 3.58 2.72 3.58
                 2.72 2.60 3.44 2.60 ;
        RECT  0.88 1.22 1.88 1.54 ;
    END
END adhalf_0

MACRO adfull_1
    CLASS CORE ;
    FOREIGN adfull_1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.64 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.42  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.66 3.96 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 2.76  LAYER metal1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.42  LAYER metal1  ;
        ANTENNAMAXAREACAR 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.82 2.98 4.50 2.98 4.50 2.46 4.38 2.34 3.04 2.34 3.04 3.04
                 2.72 3.04 2.72 2.02 4.52 2.02 4.82 2.32 ;
        END
    END b
    PIN ci
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.81  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  11.59 2.62 9.90 2.62 9.90 2.34 8.91 2.34 8.91 2.42 7.19 2.42
                 7.19 2.10 8.61 2.10 8.61 2.02 10.22 2.02 10.22 2.30 11.04 2.30
                 11.04 2.08 11.36 2.08 11.36 2.30 11.59 2.30 ;
        END
    END ci
    PIN co
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  0.50 4.54 0.18 4.54 0.18 2.40 0.16 2.40 0.16 2.08 0.18 2.08
                 0.18 1.22 0.50 1.22 ;
        END
    END co
    PIN s
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.66  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.48 3.04 16.46 3.04 16.46 4.54 16.14 4.54 16.14 1.22
                 16.46 1.22 16.46 2.72 16.48 2.72 ;
        END
    END s
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 0.90 15.56 0.90 15.56 1.54 15.24 1.54 15.24 0.90
                 7.74 0.90 7.74 1.54 7.42 1.54 7.42 0.90 5.36 0.90 5.36 1.14
                 5.04 1.14 5.04 0.90 3.96 0.90 3.96 1.54 3.64 1.54 3.64 0.90
                 1.20 0.90 1.20 1.54 0.88 1.54 0.88 0.90 0.00 0.90 0.00 -0.90
                 16.64 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 3.58 1.20 3.58
                 1.20 4.86 3.64 4.86 3.64 4.22 3.96 4.22 3.96 4.86 7.59 4.86
                 7.59 4.22 7.91 4.22 7.91 4.86 15.35 4.86 15.35 3.58 15.67 3.58
                 15.67 4.86 16.64 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  15.80 2.56 14.88 2.56 14.88 3.90 12.11 3.90 12.11 4.54
                 11.79 4.54 11.79 3.90 11.43 3.90 11.43 4.54 11.11 4.54
                 11.11 3.58 14.56 3.58 14.56 2.18 12.15 2.18 11.51 1.54
                 11.06 1.54 11.06 1.22 12.06 1.22 12.06 1.62 12.30 1.86
                 14.88 1.86 14.88 2.24 15.80 2.24 ;
        RECT  13.87 4.22 14.87 4.54 ;
        RECT  13.82 1.22 14.82 1.54 ;
        POLYGON  13.84 3.26 9.26 3.26 9.26 3.06 5.78 3.06 5.78 2.74 9.26 2.74
                 9.26 2.66 9.58 2.66 9.58 2.94 13.52 2.94 13.52 2.66 13.84 2.66 ;
        RECT  12.49 4.22 13.49 4.54 ;
        RECT  12.44 1.22 13.44 1.54 ;
        RECT  8.29 4.22 10.71 4.54 ;
        RECT  8.12 1.22 10.68 1.54 ;
        POLYGON  10.37 3.90 7.23 3.90 7.23 4.54 6.91 4.54 6.91 3.90 1.88 3.90
                 1.88 4.54 1.56 4.54 1.56 2.46 0.82 2.46 0.82 2.14 1.56 2.14
                 1.56 1.22 1.88 1.22 1.88 3.58 5.14 3.58 5.14 2.10 6.42 2.10
                 6.42 1.22 6.74 1.22 6.74 2.42 5.46 2.42 5.46 3.58 10.37 3.58 ;
        RECT  4.34 4.22 6.52 4.54 ;
        POLYGON  6.04 1.78 4.76 1.78 4.52 1.54 4.34 1.54 4.34 1.22 4.66 1.22
                 4.90 1.46 5.72 1.46 5.72 1.22 6.04 1.22 ;
        RECT  2.26 1.22 3.26 1.54 ;
        RECT  2.26 4.22 3.26 4.54 ;
    END
END adfull_1

MACRO adfull_0
    CLASS CORE ;
    FOREIGN adfull_0 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.64 BY 5.76 ;
    SYMMETRY X Y ;
    SITE CORE ;
    PIN a
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.42  LAYER metal1  ;
        PORT
        LAYER metal1 ;
        RECT  3.36 2.66 3.96 3.04 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 2.76  LAYER metal1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.42  LAYER metal1  ;
        ANTENNAMAXAREACAR 1.14  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  4.82 2.98 4.50 2.98 4.50 2.46 4.38 2.34 3.04 2.34 3.04 3.04
                 2.72 3.04 2.72 2.02 4.52 2.02 4.82 2.32 ;
        END
    END b
    PIN ci
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.83  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  11.59 2.62 9.90 2.62 9.90 2.34 8.91 2.34 8.91 2.42 7.19 2.42
                 7.19 2.10 8.61 2.10 8.61 2.02 10.22 2.02 10.22 2.30 11.04 2.30
                 11.04 2.08 11.36 2.08 11.36 2.30 11.59 2.30 ;
        END
    END ci
    PIN co
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  0.50 4.54 0.18 4.54 0.18 2.40 0.16 2.40 0.16 2.08 0.18 2.08
                 0.18 1.22 0.50 1.22 ;
        END
    END co
    PIN s
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.20  LAYER metal1  ;
        PORT
        LAYER metal1 ;
                POLYGON  16.48 3.04 16.46 3.04 16.46 4.54 16.14 4.54 16.14 1.22
                 16.46 1.22 16.46 2.72 16.48 2.72 ;
        END
    END s
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 0.90 15.62 0.90 15.62 1.54 15.30 1.54 15.30 0.90
                 7.74 0.90 7.74 1.54 7.42 1.54 7.42 0.90 5.36 0.90 5.36 1.14
                 5.04 1.14 5.04 0.90 3.96 0.90 3.96 1.54 3.64 1.54 3.64 0.90
                 1.20 0.90 1.20 1.54 0.88 1.54 0.88 0.90 0.00 0.90 0.00 -0.90
                 16.64 -0.90 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER metal1 ;
                POLYGON  16.64 6.66 0.00 6.66 0.00 4.86 0.88 4.86 0.88 4.22 1.20 4.22
                 1.20 4.86 3.64 4.86 3.64 4.22 3.96 4.22 3.96 4.86 7.54 4.86
                 7.54 4.22 7.86 4.22 7.86 4.86 15.35 4.86 15.35 4.22 15.67 4.22
                 15.67 4.86 16.64 4.86 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        POLYGON  15.80 2.56 14.88 2.56 14.88 3.90 12.06 3.90 12.06 4.54
                 11.74 4.54 11.74 3.90 11.38 3.90 11.38 4.54 11.06 4.54
                 11.06 3.58 14.56 3.58 14.56 2.18 12.15 2.18 11.51 1.54
                 11.06 1.54 11.06 1.22 12.06 1.22 12.06 1.62 12.30 1.86
                 14.88 1.86 14.88 2.24 15.80 2.24 ;
        RECT  13.82 1.22 14.82 1.54 ;
        RECT  13.82 4.22 14.82 4.54 ;
        POLYGON  13.84 3.26 9.26 3.26 9.26 3.06 5.78 3.06 5.78 2.74 9.26 2.74
                 9.26 2.66 9.58 2.66 9.58 2.94 13.52 2.94 13.52 2.66 13.84 2.66 ;
        RECT  12.44 1.22 13.44 1.54 ;
        RECT  12.44 4.22 13.44 4.54 ;
        RECT  8.12 1.22 10.68 1.54 ;
        RECT  8.24 4.22 10.66 4.54 ;
        POLYGON  10.32 3.90 7.18 3.90 7.18 4.54 6.86 4.54 6.86 3.90 1.88 3.90
                 1.88 4.54 1.56 4.54 1.56 2.46 0.82 2.46 0.82 2.14 1.56 2.14
                 1.56 1.22 1.88 1.22 1.88 3.58 5.14 3.58 5.14 2.10 6.42 2.10
                 6.42 1.22 6.74 1.22 6.74 2.42 5.46 2.42 5.46 3.58 10.32 3.58 ;
        RECT  4.34 4.22 6.47 4.54 ;
        POLYGON  6.04 1.78 4.76 1.78 4.52 1.54 4.34 1.54 4.34 1.22 4.66 1.22
                 4.90 1.46 5.72 1.46 5.72 1.22 6.04 1.22 ;
        RECT  2.26 1.22 3.26 1.54 ;
        RECT  2.26 4.22 3.26 4.54 ;
    END
END adfull_0

END LIBRARY
