#************************************************************************/
# Copyright        : (c) All Rights Reserved 
# Company          : X-FAB Semiconductor Foundries AG 
# Address          : Haarbergstr. 67,  D-99097 Erfurt, Germany 
#
# File             : D_CELLS.lef
# Description      : Layout Exchange Format
#                  
# Technology       : XC035LV
# Lib_version      : V 4.1.2  
# Last Modified by : AKT
# DATE             : Dec 14, 2004
# 
#************************************************************************/

VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
SITE core
    SYMMETRY y  ;
    CLASS core  ;
    SIZE 1.40 BY 13.00 ;
END core
#MACRO AN211X1
#    CLASS CORE ;
#    FOREIGN AN211X1 0.00 0.00  ;
#    ORIGIN 0.00 0.00 ;
#    SIZE 8.40 BY 13.00 ;
#    SYMMETRY x y r90 ;
#    SITE core ;
#    PIN Q
#        DIRECTION OUTPUT ;
#        ANTENNADIFFAREA 1.0 ;
#        PORT
#        LAYER M1M ;
#        RECT  2.80 2.45 3.50 3.65 ;
#        RECT  2.80 3.15 6.35 3.65 ;
#        RECT  5.85 2.45 6.35 10.25 ;
#        RECT  5.85 6.75 6.55 10.25 ;
#        RECT  5.85 2.45 6.60 3.15 ;
#        RECT  5.85 8.00 6.75 8.90 ;
#        END
#    END Q
#    PIN D
#        DIRECTION INPUT ;
#        ANTENNAGATEAREA 2.43 ;
#        PORT
#        LAYER M1M ;
#        RECT  4.45 4.10 5.35 5.00 ;
#        END
#    END D
#    PIN C
#        DIRECTION INPUT ;
#        ANTENNAGATEAREA 2.43 ;
#        PORT
#        LAYER M1M ;
#        RECT  3.05 4.10 3.95 5.00 ;
#        END
#    END C
#    PIN B
#        DIRECTION INPUT ;
#        ANTENNAGATEAREA 2.78 ;
#        PORT
#        LAYER M1M ;
#        RECT  1.65 5.35 2.55 6.30 ;
#        END
#    END B
#    PIN A
#        DIRECTION INPUT ;
#        ANTENNAGATEAREA 2.78 ;
#        PORT
#        LAYER M1M ;
#        RECT  0.25 5.40 1.15 6.30 ;
#        END
#    END A
#    PIN vdd!
#        DIRECTION INOUT ;
#        USE power ;
#        SHAPE ABUTMENT ;
#        PORT
#        LAYER M1M ;
#        RECT  2.15 7.75 2.85 11.00 ;
#        RECT  0.00 11.00 8.40 13.00 ;
#        END
#    END vdd!
#    PIN gnd!
#        DIRECTION INOUT ;
#        USE ground ;
#        SHAPE ABUTMENT ;
#        PORT
#        LAYER M1M ;
#        RECT  0.45 2.00 1.15 3.80 ;
#        RECT  4.35 2.00 5.05 2.70 ;
#        RECT  0.00 0.00 8.40 2.00 ;
#        END
#    END gnd!
#    OBS
#        LAYER M1M ;
#        RECT  0.80 6.75 1.50 10.55 ;
#        RECT  0.80 6.75 4.20 7.25 ;
#        RECT  3.50 6.75 4.20 10.55 ;
#    END
#END AN211X1
MACRO AN211X2
    CLASS CORE ;
    FOREIGN AN211X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  5.60 2.45 6.30 3.65 ;
        RECT  4.40 2.95 6.30 3.65 ;
        RECT  7.25 3.15 8.15 6.30 ;
        RECT  8.65 2.45 9.40 3.65 ;
        RECT  4.40 3.15 9.40 3.65 ;
        RECT  7.25 5.80 10.60 6.30 ;
        RECT  10.05 5.80 10.60 7.10 ;
        RECT  10.05 6.40 14.10 7.10 ;
        RECT  13.40 6.40 14.10 10.55 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.55 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  5.85 4.10 6.75 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.57 ;
        PORT
        LAYER M1M ;
        RECT  4.30 5.35 5.35 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.57 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.35 2.85 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.75 1.15 11.00 ;
        RECT  3.40 9.65 4.10 11.00 ;
        RECT  6.10 7.75 6.80 11.00 ;
        RECT  15.25 9.55 15.95 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.25 3.80 ;
        RECT  2.05 2.00 2.75 3.80 ;
        RECT  7.15 2.00 7.85 2.70 ;
        RECT  10.20 2.00 16.35 3.80 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.20 6.75 2.70 10.55 ;
        RECT  2.00 8.95 2.70 10.55 ;
        RECT  4.75 6.75 5.45 10.55 ;
        RECT  2.20 6.75 8.35 7.25 ;
        RECT  7.65 6.75 8.35 10.55 ;
        RECT  7.65 8.75 11.75 9.45 ;
    END
END AN211X2
MACRO AN211X4
    CLASS CORE ;
    FOREIGN AN211X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 28.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.80 3.10 13.70 3.80 ;
        RECT  14.00 2.45 14.70 3.65 ;
        RECT  8.80 3.10 14.70 3.65 ;
        RECT  17.65 2.55 18.35 3.65 ;
        RECT  20.35 2.55 21.05 3.65 ;
        RECT  8.80 3.15 21.75 3.65 ;
        RECT  21.30 3.15 21.75 9.60 ;
        RECT  21.25 3.15 21.75 5.95 ;
        RECT  21.30 5.45 22.00 9.60 ;
        RECT  21.25 4.10 22.15 5.00 ;
        RECT  21.25 5.45 24.70 5.95 ;
        RECT  24.00 5.45 24.70 9.60 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.73 ;
        PORT
        LAYER M1M ;
        RECT  19.85 4.10 20.75 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.73 ;
        PORT
        LAYER M1M ;
        RECT  17.05 4.10 17.95 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 11.13 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.35 9.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 11.13 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.35 6.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 9.60 1.15 11.00 ;
        RECT  3.30 7.75 4.00 11.00 ;
        RECT  6.00 7.75 6.70 11.00 ;
        RECT  8.70 7.75 9.40 11.00 ;
        RECT  11.40 7.75 12.10 11.00 ;
        RECT  26.85 9.60 27.55 11.00 ;
        RECT  0.00 11.00 28.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 5.65 3.80 ;
        RECT  6.45 2.00 7.15 3.80 ;
        RECT  16.30 2.00 17.00 2.70 ;
        RECT  19.00 2.00 19.70 2.70 ;
        RECT  21.70 2.00 22.40 2.70 ;
        RECT  23.25 2.00 27.55 3.80 ;
        RECT  0.00 0.00 28.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.95 6.75 2.65 10.55 ;
        RECT  4.65 6.75 5.35 10.55 ;
        RECT  7.35 6.75 8.05 10.55 ;
        RECT  10.05 6.75 10.75 10.55 ;
        RECT  1.95 6.75 13.45 7.25 ;
        RECT  12.75 6.40 13.45 10.55 ;
        RECT  14.10 5.45 14.80 9.60 ;
        RECT  15.45 6.40 16.15 10.55 ;
        RECT  16.80 5.45 17.50 9.60 ;
        RECT  18.15 6.40 18.85 10.55 ;
        RECT  12.75 10.05 18.85 10.55 ;
        RECT  14.10 5.45 20.65 5.95 ;
        RECT  19.95 5.45 20.65 10.55 ;
        RECT  22.65 6.40 23.35 10.55 ;
        RECT  25.35 6.75 26.05 10.55 ;
        RECT  19.95 10.05 26.05 10.55 ;
    END
END AN211X4
#MACRO AN21X1
#    CLASS CORE ;
#    FOREIGN AN21X1 0.00 0.00  ;
#    ORIGIN 0.00 0.00 ;
#    SIZE 7.00 BY 13.00 ;
#    SYMMETRY x y r90 ;
#    SITE core ;
#    PIN Q
#        DIRECTION OUTPUT ;
#        ANTENNADIFFAREA 1.0 ;
#        PORT
#        LAYER M1M ;
#        RECT  2.80 2.95 3.50 3.65 ;
#        RECT  3.00 2.95 3.50 4.60 ;
#        RECT  4.50 6.90 5.20 10.55 ;
#        RECT  3.00 4.10 6.75 4.60 ;
#        RECT  5.85 4.10 6.35 7.40 ;
#        RECT  4.50 6.90 6.35 7.40 ;
#        RECT  5.85 4.10 6.75 5.00 ;
#        END
#    END Q
#    PIN C
#        DIRECTION INPUT ;
#        ANTENNAGATEAREA 1.75 ;
#        PORT
#        LAYER M1M ;
#        RECT  4.45 5.40 5.35 6.30 ;
#        END
#    END C
#    PIN B
#        DIRECTION INPUT ;
#        ANTENNAGATEAREA 2.10 ;
#        PORT
#        LAYER M1M ;
#        RECT  0.25 5.40 1.15 6.30 ;
#        END
#    END B
#    PIN A
#        DIRECTION INPUT ;
#        ANTENNAGATEAREA 2.10 ;
#        PORT
#        LAYER M1M ;
#        RECT  1.65 5.40 2.95 6.30 ;
#        END
#    END A
#    PIN vdd!
#        DIRECTION INOUT ;
#        USE power ;
#        SHAPE ABUTMENT ;
#        PORT
#        LAYER M1M ;
#        RECT  1.80 7.85 2.50 11.00 ;
#        RECT  0.00 11.00 7.00 13.00 ;
#        END
#    END vdd!
#    PIN gnd!
#        DIRECTION INOUT ;
#        USE ground ;
#        SHAPE ABUTMENT ;
#        PORT
#        LAYER M1M ;
#        RECT  0.45 2.00 1.15 4.50 ;
#        RECT  4.15 2.00 4.85 3.65 ;
#        RECT  5.85 2.00 6.55 3.55 ;
#        RECT  0.00 0.00 7.00 2.00 ;
#        END
#    END gnd!
#    OBS
#        LAYER M1M ;
#        RECT  0.45 6.90 1.15 10.55 ;
#        RECT  0.45 6.90 3.85 7.40 ;
#        RECT  3.15 6.90 3.85 10.55 ;
#    END
#END AN21X1
MACRO AN21X2
    CLASS CORE ;
    FOREIGN AN21X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  5.75 2.50 6.45 4.10 ;
        RECT  5.95 2.50 6.45 4.95 ;
        RECT  5.95 4.45 9.15 4.95 ;
        RECT  8.65 4.45 9.15 9.60 ;
        RECT  8.65 5.40 9.25 9.60 ;
        RECT  8.65 7.20 9.40 9.60 ;
        RECT  8.65 5.40 9.55 6.30 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.50 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.20 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.20 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.20 1.15 11.00 ;
        RECT  3.15 7.85 3.85 11.00 ;
        RECT  5.85 7.85 6.55 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 2.05 4.70 ;
        RECT  2.90 2.00 3.60 4.50 ;
        RECT  7.10 2.00 7.80 4.00 ;
        RECT  8.60 2.00 10.75 4.00 ;
        RECT  9.60 2.00 10.75 4.70 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 6.90 2.50 10.55 ;
        RECT  4.50 6.90 5.20 10.55 ;
        RECT  1.80 6.90 8.05 7.40 ;
        RECT  7.35 6.90 8.05 10.55 ;
        RECT  10.05 7.20 10.75 10.55 ;
        RECT  7.35 10.05 10.75 10.55 ;
    END
END AN21X2
MACRO AN21X4
    CLASS CORE ;
    FOREIGN AN21X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  5.20 4.10 10.95 4.30 ;
        RECT  9.90 2.45 10.60 4.30 ;
        RECT  10.05 2.45 10.60 5.00 ;
        RECT  5.20 3.60 10.60 4.30 ;
        RECT  10.05 4.10 10.95 5.00 ;
        RECT  11.40 4.45 11.90 9.60 ;
        RECT  11.40 6.75 12.10 9.60 ;
        RECT  12.75 2.50 13.45 4.95 ;
        RECT  10.05 4.45 13.45 4.95 ;
        RECT  11.40 6.75 14.80 7.25 ;
        RECT  14.10 6.75 14.80 10.55 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 7.00 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 8.40 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 8.40 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.70 1.15 11.00 ;
        RECT  3.15 7.70 3.85 11.00 ;
        RECT  5.85 7.70 6.55 11.00 ;
        RECT  8.55 7.70 9.25 11.00 ;
        RECT  15.60 9.75 16.30 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 2.05 4.35 ;
        RECT  2.85 2.00 3.55 4.30 ;
        RECT  11.40 2.00 12.10 4.00 ;
        RECT  14.10 2.00 14.80 4.00 ;
        RECT  15.60 2.00 16.30 4.20 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 6.75 2.50 10.55 ;
        RECT  4.50 6.75 5.20 10.55 ;
        RECT  7.20 6.75 7.90 10.55 ;
        RECT  1.80 6.75 10.75 7.25 ;
        RECT  10.05 6.75 10.75 10.55 ;
        RECT  12.75 7.70 13.45 10.55 ;
        RECT  10.05 10.05 13.45 10.55 ;
    END
END AN21X4
MACRO AN221X1
    CLASS CORE ;
    FOREIGN AN221X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  3.50 3.25 9.15 3.65 ;
        RECT  3.50 2.55 4.20 3.65 ;
        RECT  7.35 3.05 8.05 3.75 ;
        RECT  3.50 3.15 8.05 3.65 ;
        RECT  7.55 6.75 8.25 10.55 ;
        RECT  7.35 3.25 9.15 3.75 ;
        RECT  8.65 3.25 9.15 7.65 ;
        RECT  8.65 6.65 9.55 7.65 ;
        RECT  7.55 6.75 9.55 7.65 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  7.15 5.35 8.15 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  5.40 4.10 6.75 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 3.95 5.00 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  1.65 4.10 2.55 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.50 7.55 4.20 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.15 2.00 1.85 3.65 ;
        RECT  5.85 2.00 6.55 2.70 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.80 5.55 1.50 10.55 ;
        RECT  2.15 6.55 2.85 10.55 ;
        RECT  2.15 6.55 5.55 7.05 ;
        RECT  4.85 6.55 5.55 10.55 ;
        RECT  0.80 5.55 6.70 6.05 ;
        RECT  6.20 5.55 6.70 10.40 ;
        RECT  6.20 7.80 6.90 10.40 ;
    END
END AN221X1
#MACRO AN221X2
#    CLASS CORE ;
#    FOREIGN AN221X2 0.00 0.00  ;
#    ORIGIN 0.00 0.00 ;
#    SIZE 18.20 BY 13.00 ;
#    SYMMETRY x y r90 ;
#    SITE core ;
#    PIN Q
#        DIRECTION OUTPUT ;
#        ANTENNADIFFAREA 1.0 ;
#        PORT
#        LAYER M1M ;
#        RECT  4.60 3.05 5.30 3.75 ;
#        RECT  5.85 2.45 6.55 3.55 ;
#        RECT  7.10 3.05 7.80 3.75 ;
#        RECT  10.95 2.85 11.90 3.55 ;
#        RECT  4.60 3.05 11.90 3.55 ;
#        RECT  11.40 2.85 11.90 5.00 ;
#        RECT  11.40 4.10 12.35 5.00 ;
#        RECT  11.40 4.50 15.05 5.00 ;
#        RECT  14.55 4.50 15.05 9.55 ;
#        RECT  14.55 7.85 15.25 9.55 ;
#        END
#    END Q
#    PIN E
#        DIRECTION INPUT ;
#        ANTENNAGATEAREA 4.90 ;
#        PORT
#        LAYER M1M ;
#        RECT  10.05 4.10 10.95 5.00 ;
#        END
#    END E
#    PIN D
#        DIRECTION INPUT ;
#        ANTENNAGATEAREA 5.58 ;
#        PORT
#        LAYER M1M ;
#        RECT  0.25 5.40 1.15 6.30 ;
#        RECT  7.50 4.25 8.00 5.95 ;
#        RECT  0.25 5.45 8.00 5.95 ;
#        RECT  7.50 4.25 8.20 4.95 ;
#        END
#    END D
#    PIN C
#        DIRECTION INPUT ;
#        ANTENNAGATEAREA 5.60 ;
#        PORT
#        LAYER M1M ;
#        RECT  8.65 4.10 9.55 5.00 ;
#        END
#    END C
#    PIN B
#        DIRECTION INPUT ;
#        ANTENNAGATEAREA 5.60 ;
#        PORT
#        LAYER M1M ;
#        RECT  5.85 4.10 6.75 5.00 ;
#        END
#    END B
#    PIN A
#        DIRECTION INPUT ;
#        ANTENNAGATEAREA 5.60 ;
#        PORT
#        LAYER M1M ;
#        RECT  2.90 4.10 3.95 5.00 ;
#        END
#    END A
#    PIN vdd!
#        DIRECTION INOUT ;
#        USE power ;
#        SHAPE ABUTMENT ;
#        PORT
#        LAYER M1M ;
#        RECT  4.90 8.30 5.60 11.00 ;
#        RECT  7.60 8.30 8.30 11.00 ;
#        RECT  0.00 11.00 18.20 13.00 ;
#        END
#    END vdd!
#    PIN gnd!
#        DIRECTION INOUT ;
#        USE ground ;
#        SHAPE ABUTMENT ;
#        PORT
#        LAYER M1M ;
#        RECT  0.45 2.00 1.40 3.80 ;
#        RECT  2.25 2.00 2.95 3.65 ;
#        RECT  9.45 2.00 10.15 2.60 ;
#        RECT  12.55 2.00 17.75 3.65 ;
#        RECT  12.70 2.00 17.75 3.80 ;
#        RECT  0.00 0.00 18.20 2.00 ;
#        END
#    END gnd!
#    OBS
#        LAYER M1M ;
#        RECT  0.85 8.10 1.55 10.55 ;
#        RECT  2.20 6.40 2.90 9.60 ;
#        RECT  3.55 7.35 4.25 10.55 ;
#        RECT  0.85 10.05 4.25 10.55 ;
#        RECT  6.25 7.35 6.95 10.55 ;
#        RECT  3.55 7.35 9.65 7.85 ;
#        RECT  8.95 7.35 9.65 10.55 ;
#        RECT  10.30 6.40 11.00 9.60 ;
#        RECT  11.65 7.35 12.35 10.55 ;
#        RECT  8.95 10.05 12.35 10.55 ;
#        RECT  2.20 6.40 13.90 6.90 ;
#        RECT  13.20 6.40 13.90 10.50 ;
#        RECT  15.90 6.95 16.60 10.50 ;
#        RECT  13.20 10.00 16.60 10.50 ;
#    END
#END AN221X2
MACRO AN221X4
    CLASS CORE ;
    FOREIGN AN221X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 33.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  13.10 2.45 13.80 3.80 ;
        RECT  8.55 3.10 18.05 3.80 ;
        RECT  22.15 2.50 22.85 3.65 ;
        RECT  8.55 3.15 22.85 3.65 ;
        RECT  22.35 2.50 22.85 5.95 ;
        RECT  22.35 5.45 27.75 5.95 ;
        RECT  26.90 5.40 27.60 9.60 ;
        RECT  26.85 5.40 27.75 6.30 ;
        RECT  26.85 5.40 30.30 5.90 ;
        RECT  22.35 5.45 30.30 5.90 ;
        RECT  29.60 5.40 30.30 9.60 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.73 ;
        PORT
        LAYER M1M ;
        RECT  25.45 4.10 26.35 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 11.13 ;
        PORT
        LAYER M1M ;
        RECT  18.45 4.10 19.35 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 11.13 ;
        PORT
        LAYER M1M ;
        RECT  19.85 4.10 20.75 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 11.13 ;
        PORT
        LAYER M1M ;
        RECT  7.25 4.10 8.15 5.00 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 11.13 ;
        PORT
        LAYER M1M ;
        RECT  5.85 4.10 6.75 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 9.60 1.20 11.00 ;
        RECT  2.15 7.35 2.85 11.00 ;
        RECT  4.85 7.35 5.55 11.00 ;
        RECT  7.55 7.35 8.25 11.00 ;
        RECT  10.25 7.35 10.95 11.00 ;
        RECT  12.95 7.35 13.65 11.00 ;
        RECT  32.45 9.60 33.15 11.00 ;
        RECT  0.00 11.00 33.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 4.75 3.80 ;
        RECT  5.55 2.00 6.25 3.60 ;
        RECT  20.65 2.00 21.35 2.70 ;
        RECT  23.50 2.00 24.20 3.60 ;
        RECT  25.25 2.00 33.15 2.95 ;
        RECT  27.05 2.00 33.15 3.80 ;
        RECT  0.00 0.00 33.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.50 6.40 4.20 10.55 ;
        RECT  6.20 6.40 6.90 10.55 ;
        RECT  8.90 6.40 9.60 10.55 ;
        RECT  11.60 6.40 12.30 9.80 ;
        RECT  14.75 7.35 15.45 10.55 ;
        RECT  16.10 6.40 16.80 9.60 ;
        RECT  17.45 7.35 18.15 10.55 ;
        RECT  18.80 6.40 19.50 9.60 ;
        RECT  20.15 7.35 20.85 10.55 ;
        RECT  21.50 6.40 22.20 9.60 ;
        RECT  22.85 7.35 23.55 10.55 ;
        RECT  3.50 6.40 24.90 6.90 ;
        RECT  24.20 6.40 24.90 9.60 ;
        RECT  25.55 6.40 26.25 10.55 ;
        RECT  28.25 6.40 28.95 10.55 ;
        RECT  30.95 6.60 31.65 10.55 ;
        RECT  14.75 10.05 31.65 10.55 ;
    END
END AN221X4
MACRO AN222X1
    CLASS CORE ;
    FOREIGN AN222X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  3.60 2.65 4.30 3.65 ;
        RECT  7.55 5.80 8.25 9.60 ;
        RECT  9.20 2.65 9.90 3.65 ;
        RECT  3.60 3.15 10.55 3.65 ;
        RECT  10.05 3.15 10.55 6.30 ;
        RECT  10.05 5.40 10.95 6.30 ;
        RECT  7.55 5.80 10.95 6.30 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.55 5.00 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  7.25 4.10 8.15 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  5.50 4.10 6.75 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 3.95 5.00 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  1.65 4.10 2.55 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.50 7.40 4.20 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.25 2.00 1.95 3.65 ;
        RECT  5.95 2.00 7.55 2.70 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.80 5.45 1.50 10.55 ;
        RECT  2.15 6.45 2.85 10.55 ;
        RECT  2.15 6.45 5.55 6.95 ;
        RECT  4.85 6.45 5.55 10.55 ;
        RECT  0.80 5.45 6.90 5.95 ;
        RECT  6.20 5.45 6.90 10.55 ;
        RECT  8.90 7.00 9.60 10.55 ;
        RECT  6.20 10.05 9.60 10.55 ;
    END
END AN222X1
MACRO AN222X2
    CLASS CORE ;
    FOREIGN AN222X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.60 3.05 5.30 3.75 ;
        RECT  5.85 2.45 6.55 3.55 ;
        RECT  7.10 3.05 7.80 3.75 ;
        RECT  4.60 3.05 10.75 3.55 ;
        RECT  10.25 3.05 10.75 5.00 ;
        RECT  14.25 2.45 14.55 5.00 ;
        RECT  13.85 2.45 14.55 3.65 ;
        RECT  14.25 2.95 15.15 5.00 ;
        RECT  10.25 4.50 15.15 5.00 ;
        RECT  14.65 2.95 15.15 5.95 ;
        RECT  13.85 2.95 15.80 3.65 ;
        RECT  15.40 5.45 16.10 9.60 ;
        RECT  14.65 5.45 18.80 5.95 ;
        RECT  18.10 5.45 18.80 9.60 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.60 ;
        PORT
        LAYER M1M ;
        RECT  15.65 4.10 16.55 5.00 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.58 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.58 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        RECT  7.50 4.25 8.00 5.95 ;
        RECT  0.25 5.45 8.00 5.95 ;
        RECT  7.50 4.25 8.20 4.95 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.60 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.55 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.60 ;
        PORT
        LAYER M1M ;
        RECT  5.85 4.10 6.75 5.00 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.60 ;
        PORT
        LAYER M1M ;
        RECT  2.90 4.10 3.95 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  4.90 8.30 5.60 11.00 ;
        RECT  7.60 8.30 8.30 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.60 2.00 1.30 3.80 ;
        RECT  2.25 2.00 2.95 3.65 ;
        RECT  9.45 2.00 10.15 2.60 ;
        RECT  11.20 2.00 12.80 3.80 ;
        RECT  17.45 2.00 18.15 3.65 ;
        RECT  18.95 2.00 20.55 3.80 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.85 8.10 1.55 10.55 ;
        RECT  2.20 6.40 2.90 9.60 ;
        RECT  3.55 7.35 4.25 10.55 ;
        RECT  0.85 10.05 4.25 10.55 ;
        RECT  6.25 7.35 6.95 10.55 ;
        RECT  3.55 7.35 9.65 7.85 ;
        RECT  8.95 7.35 9.65 10.55 ;
        RECT  10.30 6.40 11.00 9.60 ;
        RECT  11.65 7.35 12.35 10.55 ;
        RECT  8.95 10.05 12.35 10.55 ;
        RECT  2.20 6.40 14.75 6.90 ;
        RECT  14.05 6.40 14.75 10.55 ;
        RECT  16.75 6.50 17.45 10.55 ;
        RECT  19.45 8.10 20.15 10.55 ;
        RECT  14.05 10.05 20.15 10.55 ;
    END
END AN222X2
MACRO AN222X4
    CLASS CORE ;
    FOREIGN AN222X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 39.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  13.10 2.45 13.80 3.80 ;
        RECT  8.55 3.10 18.05 3.80 ;
        RECT  25.45 2.45 26.15 3.60 ;
        RECT  8.55 3.10 30.70 3.60 ;
        RECT  26.90 3.10 27.35 9.60 ;
        RECT  26.85 3.10 27.35 6.30 ;
        RECT  26.90 5.40 27.60 9.60 ;
        RECT  26.85 5.40 27.75 6.30 ;
        RECT  29.60 5.45 30.30 9.60 ;
        RECT  26.35 3.10 30.70 3.80 ;
        RECT  32.30 5.45 33.00 9.60 ;
        RECT  26.85 5.45 35.70 5.95 ;
        RECT  35.00 5.45 35.70 9.60 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 11.13 ;
        PORT
        LAYER M1M ;
        RECT  31.05 4.10 31.95 5.00 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 11.13 ;
        PORT
        LAYER M1M ;
        RECT  32.45 4.10 33.35 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 11.13 ;
        PORT
        LAYER M1M ;
        RECT  18.45 4.05 19.35 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 11.13 ;
        PORT
        LAYER M1M ;
        RECT  19.85 4.10 20.75 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 11.13 ;
        PORT
        LAYER M1M ;
        RECT  7.25 4.10 8.15 5.00 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 11.13 ;
        PORT
        LAYER M1M ;
        RECT  5.85 4.10 6.75 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 9.60 1.20 11.00 ;
        RECT  2.15 7.35 2.85 11.00 ;
        RECT  4.85 7.35 5.55 11.00 ;
        RECT  7.55 7.35 8.25 11.00 ;
        RECT  10.25 7.35 10.95 11.00 ;
        RECT  12.95 7.35 13.65 11.00 ;
        RECT  37.95 9.60 38.65 11.00 ;
        RECT  0.00 11.00 39.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 4.75 3.80 ;
        RECT  5.55 2.00 6.25 3.60 ;
        RECT  20.65 2.00 21.35 2.65 ;
        RECT  33.00 2.00 33.70 3.60 ;
        RECT  34.50 2.00 38.75 3.80 ;
        RECT  0.00 0.00 39.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.50 6.40 4.20 10.55 ;
        RECT  6.20 6.40 6.90 10.55 ;
        RECT  8.90 6.40 9.60 10.55 ;
        RECT  11.60 6.40 12.30 9.80 ;
        RECT  14.75 7.35 15.45 10.55 ;
        RECT  16.10 6.40 16.80 9.60 ;
        RECT  17.45 7.35 18.15 10.55 ;
        RECT  18.80 6.40 19.50 9.60 ;
        RECT  20.15 7.35 20.85 10.55 ;
        RECT  21.50 6.40 22.20 9.60 ;
        RECT  22.85 7.35 23.55 10.55 ;
        RECT  3.50 6.40 24.90 6.90 ;
        RECT  24.20 6.40 24.90 9.60 ;
        RECT  25.55 6.40 26.25 10.55 ;
        RECT  28.25 6.40 28.95 10.55 ;
        RECT  30.95 6.40 31.65 10.55 ;
        RECT  33.65 6.40 34.35 10.55 ;
        RECT  36.35 6.75 37.05 10.55 ;
        RECT  14.75 10.05 37.05 10.55 ;
    END
END AN222X4
MACRO AN22X1
    CLASS CORE ;
    FOREIGN AN22X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.65 4.45 2.15 9.60 ;
        RECT  1.65 7.45 2.55 9.60 ;
        RECT  3.15 2.45 3.85 4.95 ;
        RECT  1.65 4.45 3.85 4.95 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  2.75 5.40 3.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  4.40 5.35 5.35 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  4.50 7.85 5.20 11.00 ;
        RECT  0.00 11.00 7.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.80 2.00 1.50 4.00 ;
        RECT  5.50 2.00 6.20 4.00 ;
        RECT  0.00 0.00 7.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 7.20 1.15 10.55 ;
        RECT  3.15 6.90 3.85 10.55 ;
        RECT  0.45 10.05 3.85 10.55 ;
        RECT  3.15 6.90 6.55 7.40 ;
        RECT  5.85 6.90 6.55 10.55 ;
    END
END AN22X1
MACRO AN22X2
    CLASS CORE ;
    FOREIGN AN22X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.50 6.90 1.20 10.55 ;
        RECT  3.20 6.90 3.90 9.60 ;
        RECT  5.85 3.80 6.75 7.40 ;
        RECT  0.50 6.90 6.75 7.40 ;
        RECT  6.20 2.45 6.75 9.60 ;
        RECT  5.90 3.80 6.75 9.60 ;
        RECT  6.20 2.45 6.90 4.50 ;
        RECT  5.70 3.80 7.40 4.50 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.20 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.20 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.35 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.20 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.35 12.35 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.20 ;
        PORT
        LAYER M1M ;
        RECT  7.20 5.35 8.15 6.35 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  8.75 7.85 9.45 11.00 ;
        RECT  11.45 7.85 12.15 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 2.55 4.70 ;
        RECT  3.35 2.00 4.05 4.50 ;
        RECT  9.05 2.00 9.75 4.50 ;
        RECT  10.55 2.00 13.55 4.70 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.85 7.85 2.55 10.55 ;
        RECT  4.55 7.85 5.25 10.55 ;
        RECT  7.40 6.90 8.10 10.55 ;
        RECT  1.85 10.05 8.10 10.55 ;
        RECT  10.10 6.90 10.80 10.55 ;
        RECT  7.40 6.90 13.50 7.40 ;
        RECT  12.80 6.90 13.50 10.55 ;
    END
END AN22X2
MACRO AN22X4
    CLASS CORE ;
    FOREIGN AN22X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.15 2.45 10.85 4.30 ;
        RECT  12.85 3.60 13.75 5.00 ;
        RECT  13.25 3.60 13.75 9.60 ;
        RECT  13.10 6.75 13.80 9.60 ;
        RECT  5.20 3.60 15.80 4.30 ;
        RECT  15.80 6.75 16.50 9.60 ;
        RECT  13.10 6.75 19.20 7.25 ;
        RECT  18.50 6.75 19.20 9.60 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 8.40 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 8.40 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 8.40 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 8.40 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.70 1.15 11.00 ;
        RECT  3.15 7.70 3.85 11.00 ;
        RECT  5.85 7.70 6.55 11.00 ;
        RECT  8.55 7.70 9.25 11.00 ;
        RECT  10.15 7.70 10.85 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 2.05 4.35 ;
        RECT  2.85 2.00 3.55 4.30 ;
        RECT  17.45 2.00 18.15 4.30 ;
        RECT  18.95 2.00 20.55 4.30 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 6.75 2.50 10.55 ;
        RECT  4.50 6.75 5.20 10.55 ;
        RECT  7.20 6.75 7.90 10.55 ;
        RECT  1.80 6.75 12.45 7.25 ;
        RECT  11.75 6.75 12.45 10.55 ;
        RECT  14.45 7.70 15.15 10.55 ;
        RECT  17.15 7.70 17.85 10.55 ;
        RECT  19.85 7.15 20.55 10.55 ;
        RECT  11.75 10.05 20.55 10.55 ;
    END
END AN22X4
MACRO AN311X1
    CLASS CORE ;
    FOREIGN AN311X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  3.80 2.45 4.50 3.65 ;
        RECT  6.80 2.55 7.70 3.65 ;
        RECT  3.80 3.15 7.70 3.65 ;
        RECT  7.20 2.55 7.70 10.40 ;
        RECT  7.20 6.65 7.90 10.40 ;
        RECT  7.20 8.00 8.15 8.90 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  5.85 4.10 6.75 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  4.45 4.10 5.40 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 3.95 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.35 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.80 8.10 1.50 11.00 ;
        RECT  3.50 7.70 4.20 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.65 ;
        RECT  5.30 2.00 6.00 2.70 ;
        RECT  8.55 2.00 9.25 3.80 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.15 6.75 2.85 10.55 ;
        RECT  2.15 6.75 5.55 7.25 ;
        RECT  4.85 6.75 5.55 10.55 ;
    END
END AN311X1
MACRO AN311X2
    CLASS CORE ;
    FOREIGN AN311X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  7.90 2.45 8.60 4.80 ;
        RECT  5.55 4.10 8.60 4.80 ;
        RECT  14.20 2.45 15.15 3.60 ;
        RECT  7.90 3.10 15.15 3.60 ;
        RECT  14.45 2.45 14.95 6.25 ;
        RECT  14.25 2.45 15.15 3.70 ;
        RECT  14.45 5.75 16.25 6.25 ;
        RECT  15.55 5.75 16.25 7.80 ;
        RECT  15.55 7.10 19.15 7.80 ;
        RECT  18.45 7.10 19.15 10.55 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  15.65 4.10 16.55 5.00 ;
        RECT  15.40 4.30 16.55 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  12.85 4.10 13.75 5.00 ;
        RECT  12.85 4.30 14.00 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.35 3.95 6.30 ;
        RECT  3.05 5.60 4.25 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.35 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.40 1.15 11.00 ;
        RECT  0.45 10.40 2.60 11.00 ;
        RECT  4.20 7.70 4.90 11.00 ;
        RECT  2.80 7.70 6.30 8.40 ;
        RECT  7.95 7.70 8.65 11.00 ;
        RECT  6.55 10.40 10.05 11.00 ;
        RECT  10.30 7.70 12.40 8.40 ;
        RECT  11.70 7.70 12.40 11.00 ;
        RECT  0.00 11.00 19.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.25 3.80 ;
        RECT  2.05 2.00 2.75 4.50 ;
        RECT  9.40 2.00 12.05 2.65 ;
        RECT  12.85 2.00 13.55 2.65 ;
        RECT  15.60 2.00 16.30 3.15 ;
        RECT  17.10 2.00 19.15 3.75 ;
        RECT  0.00 0.00 19.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 6.75 2.30 9.75 ;
        RECT  1.80 9.05 3.55 9.75 ;
        RECT  6.80 6.75 7.30 9.75 ;
        RECT  5.55 9.05 7.30 9.75 ;
        RECT  9.30 6.75 9.80 9.75 ;
        RECT  9.30 9.05 11.05 9.75 ;
        RECT  1.80 6.75 13.90 7.25 ;
        RECT  13.20 5.75 13.90 10.15 ;
        RECT  13.20 9.45 16.80 10.15 ;
    END
END AN311X2
MACRO AN311X4
    CLASS CORE ;
    FOREIGN AN311X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 36.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  21.85 2.45 22.55 4.85 ;
        RECT  13.55 4.10 22.55 4.85 ;
        RECT  26.20 2.45 26.70 4.85 ;
        RECT  26.20 2.45 26.90 3.15 ;
        RECT  28.25 4.10 29.20 5.00 ;
        RECT  28.90 2.45 29.20 9.60 ;
        RECT  28.70 4.10 29.20 7.25 ;
        RECT  28.90 2.45 29.40 4.85 ;
        RECT  13.55 4.35 29.40 4.85 ;
        RECT  28.80 6.75 29.50 9.60 ;
        RECT  28.90 2.45 29.60 3.15 ;
        RECT  31.50 6.75 32.20 9.60 ;
        RECT  28.70 6.75 34.90 7.25 ;
        RECT  34.20 6.75 34.90 10.55 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  29.65 5.35 30.55 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  26.75 5.40 27.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.40 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.10 1.15 11.00 ;
        RECT  3.15 6.50 3.85 11.00 ;
        RECT  5.85 6.50 6.55 11.00 ;
        RECT  8.55 7.80 9.25 11.00 ;
        RECT  11.25 7.80 11.95 11.00 ;
        RECT  13.95 7.80 14.65 11.00 ;
        RECT  16.65 7.80 17.35 11.00 ;
        RECT  19.35 7.80 20.05 11.00 ;
        RECT  0.00 11.00 36.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 9.25 3.80 ;
        RECT  10.05 2.00 10.75 4.15 ;
        RECT  23.35 2.00 24.05 3.80 ;
        RECT  24.85 2.00 25.55 3.65 ;
        RECT  27.55 2.00 28.25 3.65 ;
        RECT  30.25 2.00 30.95 3.65 ;
        RECT  31.75 2.00 35.90 3.80 ;
        RECT  0.00 0.00 36.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 5.55 2.50 10.55 ;
        RECT  4.50 5.55 5.20 10.55 ;
        RECT  1.80 5.55 7.90 6.05 ;
        RECT  7.20 5.55 7.90 10.55 ;
        RECT  9.90 6.85 10.60 10.55 ;
        RECT  12.60 6.85 13.30 10.55 ;
        RECT  15.30 6.85 16.00 10.55 ;
        RECT  18.00 6.85 18.70 10.55 ;
        RECT  7.20 6.85 21.40 7.35 ;
        RECT  20.70 6.85 21.40 10.55 ;
        RECT  22.05 6.85 22.75 9.60 ;
        RECT  23.40 7.90 24.10 10.55 ;
        RECT  24.75 6.85 25.45 9.60 ;
        RECT  26.10 7.90 26.80 10.55 ;
        RECT  20.70 10.05 26.80 10.55 ;
        RECT  22.05 6.85 28.15 7.35 ;
        RECT  27.45 6.85 28.15 10.55 ;
        RECT  30.15 7.70 30.85 10.55 ;
        RECT  32.85 7.70 33.55 10.55 ;
        RECT  27.45 10.05 33.55 10.55 ;
    END
END AN311X4
MACRO AN31X1
    CLASS CORE ;
    FOREIGN AN31X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  3.80 2.60 4.50 4.90 ;
        RECT  3.80 4.40 6.35 4.90 ;
        RECT  5.85 4.40 6.35 10.55 ;
        RECT  5.85 7.20 6.55 10.55 ;
        RECT  5.85 8.00 6.75 8.90 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.40 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.35 3.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.35 2.60 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.20 1.15 11.00 ;
        RECT  3.15 7.85 3.85 11.00 ;
        RECT  0.00 11.00 7.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 4.20 ;
        RECT  5.30 2.00 6.00 3.70 ;
        RECT  0.00 0.00 7.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 6.90 2.50 10.55 ;
        RECT  1.80 6.90 5.20 7.40 ;
        RECT  4.50 6.90 5.20 10.55 ;
    END
END AN31X1
MACRO AN31X2
    CLASS CORE ;
    FOREIGN AN31X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.45 2.45 9.15 4.55 ;
        RECT  6.10 3.85 9.15 4.55 ;
        RECT  8.65 2.45 9.15 6.30 ;
        RECT  8.65 5.40 9.55 6.30 ;
        RECT  8.65 5.80 10.45 6.30 ;
        RECT  9.95 5.80 10.45 9.60 ;
        RECT  9.95 7.15 10.65 9.60 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.50 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.35 8.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.35 5.35 6.40 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 7.85 2.55 11.00 ;
        RECT  4.55 7.85 5.25 11.00 ;
        RECT  7.25 7.85 7.95 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.75 4.50 ;
        RECT  2.55 2.00 3.25 4.50 ;
        RECT  9.80 2.00 10.50 4.25 ;
        RECT  11.40 2.00 12.10 4.70 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.50 6.90 1.20 10.55 ;
        RECT  3.20 6.90 3.90 10.55 ;
        RECT  5.90 6.90 6.60 10.55 ;
        RECT  0.50 6.90 9.30 7.40 ;
        RECT  8.60 6.90 9.30 10.55 ;
        RECT  11.30 7.15 12.00 10.55 ;
        RECT  8.60 10.05 12.00 10.55 ;
    END
END AN31X2
#MACRO AN31X4
#    CLASS CORE ;
#    FOREIGN AN31X4 0.00 0.00  ;
#    ORIGIN 0.00 0.00 ;
#    SIZE 23.80 BY 13.00 ;
#    SYMMETRY x y r90 ;
#    SITE core ;
#    PIN Q
#        DIRECTION OUTPUT ;
#        ANTENNADIFFAREA 1.0 ;
#        PORT
#        LAYER M1M ;
#        RECT  18.45 4.10 19.35 6.30 ;
#        RECT  18.90 2.45 19.30 9.60 ;
#        RECT  18.60 4.10 19.30 9.60 ;
#        RECT  18.90 2.45 19.35 7.25 ;
#        RECT  18.60 4.10 19.35 7.25 ;
#        RECT  18.90 2.45 19.60 4.80 ;
#        RECT  10.55 4.10 19.60 4.80 ;
#        RECT  18.60 6.75 22.00 7.25 ;
#        RECT  21.30 6.75 22.00 9.60 ;
#        END
#    END Q
#    PIN D
#        DIRECTION INPUT ;
#        ANTENNAGATEAREA 7.00 ;
#        PORT
#        LAYER M1M ;
#        RECT  19.85 5.40 20.75 6.30 ;
#        END
#    END D
#    PIN C
#        DIRECTION INPUT ;
#        ANTENNAGATEAREA 9.80 ;
#        PORT
#        LAYER M1M ;
#        RECT  12.85 5.35 13.75 6.30 ;
#        END
#    END C
#    PIN B
#        DIRECTION INPUT ;
#        ANTENNAGATEAREA 9.80 ;
#        PORT
#        LAYER M1M ;
#        RECT  8.65 5.35 9.55 6.30 ;
#        END
#    END B
#    PIN A
#        DIRECTION INPUT ;
#        ANTENNAGATEAREA 9.80 ;
#        PORT
#        LAYER M1M ;
#        RECT  5.85 5.40 6.75 6.30 ;
#        END
#    END A
#    PIN vdd!
#        DIRECTION INOUT ;
#        USE power ;
#        SHAPE ABUTMENT ;
#        PORT
#        LAYER M1M ;
#        RECT  2.40 7.70 3.10 11.00 ;
#        RECT  5.10 7.70 5.80 11.00 ;
#        RECT  7.80 7.70 8.50 11.00 ;
#        RECT  10.50 7.70 11.20 11.00 ;
#        RECT  13.20 7.70 13.90 11.00 ;
#        RECT  15.90 7.70 16.60 11.00 ;
#        RECT  0.00 11.00 23.80 13.00 ;
#        END
#    END vdd!
#    PIN gnd!
#        DIRECTION INOUT ;
#        USE ground ;
#        SHAPE ABUTMENT ;
#        PORT
#        LAYER M1M ;
#        RECT  0.45 2.00 6.10 4.50 ;
#        RECT  7.05 2.00 7.75 4.40 ;
#        RECT  20.25 2.00 20.95 4.60 ;
#        RECT  21.75 2.00 23.35 4.70 ;
#        RECT  0.00 0.00 23.80 2.00 ;
#        END
#    END gnd!
#    OBS
#        LAYER M1M ;
#        RECT  1.05 6.75 1.75 10.55 ;
#        RECT  3.75 6.75 4.45 10.55 ;
#        RECT  6.45 6.75 7.15 10.55 ;
#        RECT  9.15 6.75 9.85 10.55 ;
#        RECT  11.85 6.75 12.55 10.55 ;
#        RECT  14.55 6.75 15.25 10.55 ;
#        RECT  1.05 6.75 17.95 7.25 ;
#        RECT  17.25 6.75 17.95 10.55 ;
#        RECT  19.95 7.70 20.65 10.55 ;
#        RECT  22.65 7.70 23.35 10.55 ;
#        RECT  17.25 10.05 23.35 10.55 ;
#    END
#END AN31X4
MACRO AN321X1
    CLASS CORE ;
    FOREIGN AN321X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.45 4.30 11.25 4.80 ;
        RECT  5.80 2.45 6.30 3.65 ;
        RECT  3.80 2.45 6.30 3.15 ;
        RECT  9.45 2.80 10.95 3.65 ;
        RECT  5.80 3.15 10.95 3.65 ;
        RECT  10.05 2.80 10.95 3.70 ;
        RECT  10.75 2.80 10.95 10.55 ;
        RECT  10.45 2.80 10.95 4.80 ;
        RECT  10.75 4.30 11.25 10.55 ;
        RECT  10.75 7.10 11.45 10.55 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.55 5.00 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  5.85 4.10 6.75 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  7.25 4.10 8.15 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 3.95 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  1.65 4.10 2.55 5.65 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.80 8.20 1.50 11.00 ;
        RECT  3.50 7.05 4.20 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.80 ;
        RECT  7.95 2.00 8.65 2.70 ;
        RECT  11.45 2.00 12.15 3.80 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.15 6.10 2.85 10.55 ;
        RECT  2.15 6.10 5.55 6.60 ;
        RECT  4.85 6.10 5.55 10.55 ;
        RECT  6.20 6.10 6.90 9.60 ;
        RECT  7.55 7.05 8.25 10.55 ;
        RECT  4.85 10.05 8.25 10.55 ;
        RECT  6.20 6.10 10.10 6.60 ;
        RECT  9.40 6.10 10.10 10.10 ;
    END
END AN321X1
MACRO AN321X2
    CLASS CORE ;
    FOREIGN AN321X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  19.85 4.10 20.75 5.00 ;
        RECT  7.90 2.45 8.60 4.80 ;
        RECT  5.55 4.10 8.60 4.80 ;
        RECT  14.30 2.45 15.00 3.65 ;
        RECT  14.30 3.10 16.20 3.65 ;
        RECT  15.50 3.10 16.20 3.80 ;
        RECT  7.90 3.15 20.35 3.65 ;
        RECT  19.85 2.45 19.90 5.00 ;
        RECT  19.20 2.45 19.90 3.65 ;
        RECT  20.20 3.15 20.35 9.60 ;
        RECT  19.85 3.15 20.35 5.00 ;
        RECT  20.20 4.10 20.75 9.60 ;
        RECT  20.20 7.10 20.90 9.60 ;
        RECT  20.20 8.90 21.10 9.60 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.87 ;
        PORT
        LAYER M1M ;
        RECT  18.45 4.10 19.35 5.00 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.57 ;
        PORT
        LAYER M1M ;
        RECT  14.20 4.10 15.15 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.57 ;
        PORT
        LAYER M1M ;
        RECT  17.05 4.10 17.95 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.35 3.95 6.30 ;
        RECT  3.05 5.60 4.25 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.35 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.40 1.15 11.00 ;
        RECT  1.85 10.40 2.55 11.00 ;
        RECT  4.20 7.70 4.90 11.00 ;
        RECT  2.80 7.70 6.30 8.40 ;
        RECT  7.95 7.70 8.65 11.00 ;
        RECT  6.55 10.40 10.05 11.00 ;
        RECT  10.30 7.70 12.40 8.40 ;
        RECT  11.70 7.70 12.40 11.00 ;
        RECT  0.00 11.00 23.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.25 3.80 ;
        RECT  2.05 2.00 2.75 4.50 ;
        RECT  9.50 2.00 13.50 2.65 ;
        RECT  17.85 2.00 18.55 2.70 ;
        RECT  20.80 2.00 23.35 3.65 ;
        RECT  21.10 2.00 23.35 3.80 ;
        RECT  0.00 0.00 23.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 6.75 2.30 9.75 ;
        RECT  1.80 9.05 3.55 9.75 ;
        RECT  6.80 6.75 7.30 9.75 ;
        RECT  5.55 9.05 7.30 9.75 ;
        RECT  9.30 6.75 9.80 9.75 ;
        RECT  9.30 9.05 11.05 9.75 ;
        RECT  12.35 6.20 12.85 7.25 ;
        RECT  1.80 6.75 12.85 7.25 ;
        RECT  13.30 7.15 14.00 10.55 ;
        RECT  12.35 6.20 15.35 6.70 ;
        RECT  12.35 6.40 18.05 6.70 ;
        RECT  14.65 6.20 15.35 9.25 ;
        RECT  16.00 7.35 16.70 10.55 ;
        RECT  14.65 6.40 18.05 6.90 ;
        RECT  17.35 6.40 18.05 9.60 ;
        RECT  18.70 6.40 19.40 10.55 ;
        RECT  21.95 7.15 22.65 10.55 ;
        RECT  13.30 10.05 22.65 10.55 ;
    END
END AN321X2
MACRO AN321X4
    CLASS CORE ;
    FOREIGN AN321X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 44.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  21.85 2.45 22.55 4.80 ;
        RECT  13.55 4.10 22.55 4.80 ;
        RECT  31.50 3.10 32.00 4.80 ;
        RECT  13.55 4.30 32.00 4.80 ;
        RECT  31.50 3.10 38.55 3.60 ;
        RECT  33.70 3.10 38.55 3.80 ;
        RECT  36.65 5.40 37.55 6.30 ;
        RECT  37.05 3.10 37.55 9.60 ;
        RECT  37.05 6.85 37.75 9.60 ;
        RECT  37.85 2.45 38.55 4.25 ;
        RECT  37.05 3.10 38.55 4.25 ;
        RECT  39.75 6.85 40.45 9.60 ;
        RECT  37.05 6.85 43.15 7.35 ;
        RECT  42.45 6.85 43.15 10.20 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  38.05 5.40 38.95 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 11.20 ;
        PORT
        LAYER M1M ;
        RECT  32.45 4.10 33.35 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 11.20 ;
        PORT
        LAYER M1M ;
        RECT  26.85 5.35 27.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.40 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.10 1.15 11.00 ;
        RECT  3.15 6.50 3.85 11.00 ;
        RECT  5.85 6.50 6.55 11.00 ;
        RECT  8.55 7.80 9.25 11.00 ;
        RECT  11.25 7.80 11.95 11.00 ;
        RECT  13.95 7.80 14.65 11.00 ;
        RECT  16.65 7.80 17.35 11.00 ;
        RECT  19.35 7.80 20.05 11.00 ;
        RECT  0.00 11.00 44.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 9.25 3.80 ;
        RECT  10.05 2.00 10.75 4.15 ;
        RECT  23.35 2.00 29.50 3.80 ;
        RECT  30.30 2.00 31.00 3.80 ;
        RECT  39.20 2.00 39.90 4.55 ;
        RECT  40.70 2.00 44.35 4.70 ;
        RECT  0.00 0.00 44.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 5.55 2.50 10.55 ;
        RECT  4.50 5.55 5.20 10.55 ;
        RECT  1.80 5.55 7.90 6.05 ;
        RECT  7.20 5.55 7.90 10.55 ;
        RECT  9.90 6.85 10.60 10.55 ;
        RECT  12.60 6.85 13.30 10.55 ;
        RECT  15.30 6.85 16.00 10.55 ;
        RECT  18.00 6.85 18.70 10.55 ;
        RECT  7.20 6.85 21.40 7.35 ;
        RECT  20.70 6.85 21.40 10.55 ;
        RECT  22.05 6.85 22.75 9.60 ;
        RECT  23.40 7.85 24.10 10.55 ;
        RECT  24.75 6.85 25.45 9.60 ;
        RECT  26.10 7.85 26.80 10.55 ;
        RECT  27.45 6.85 28.15 9.60 ;
        RECT  28.80 7.85 29.50 10.55 ;
        RECT  30.15 6.85 30.85 9.60 ;
        RECT  31.50 7.85 32.20 10.55 ;
        RECT  32.85 6.85 33.55 9.60 ;
        RECT  34.20 7.90 34.90 10.55 ;
        RECT  20.70 10.05 34.90 10.55 ;
        RECT  22.05 6.85 36.40 7.35 ;
        RECT  35.70 6.85 36.40 10.55 ;
        RECT  38.40 7.90 39.10 10.55 ;
        RECT  41.10 7.90 41.80 10.55 ;
        RECT  35.70 10.05 41.80 10.55 ;
    END
END AN321X4
MACRO AN322X1
    CLASS CORE ;
    FOREIGN AN322X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  3.80 3.15 10.95 3.25 ;
        RECT  4.90 2.55 5.40 3.65 ;
        RECT  3.80 2.55 5.40 3.25 ;
        RECT  4.90 3.15 10.95 3.65 ;
        RECT  10.05 2.45 10.95 3.70 ;
        RECT  10.40 2.45 10.95 9.25 ;
        RECT  10.05 2.45 11.00 3.20 ;
        RECT  3.80 3.15 11.00 3.20 ;
        RECT  10.40 7.65 11.10 9.25 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  11.40 5.00 12.40 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  8.60 4.10 9.55 5.00 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  4.45 4.10 5.70 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  7.25 4.10 8.15 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 3.95 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  1.65 4.10 2.55 5.65 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.80 8.20 1.50 11.00 ;
        RECT  3.50 7.05 4.20 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.80 ;
        RECT  7.05 2.00 8.65 2.70 ;
        RECT  11.95 2.00 13.55 3.80 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.15 6.10 2.85 10.55 ;
        RECT  2.15 6.10 5.55 6.60 ;
        RECT  4.85 6.10 5.55 10.55 ;
        RECT  6.20 6.00 6.90 9.60 ;
        RECT  7.55 6.95 8.25 10.55 ;
        RECT  4.85 10.05 8.25 10.55 ;
        RECT  6.20 6.00 9.75 6.50 ;
        RECT  9.05 6.00 9.75 10.55 ;
        RECT  11.75 7.00 12.45 10.55 ;
        RECT  9.05 10.05 12.45 10.55 ;
    END
END AN322X1
MACRO AN322X2
    CLASS CORE ;
    FOREIGN AN322X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 26.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  7.90 2.45 8.60 4.80 ;
        RECT  5.55 4.10 8.60 4.80 ;
        RECT  14.30 2.45 15.00 3.65 ;
        RECT  14.30 3.10 16.20 3.65 ;
        RECT  15.50 3.10 16.20 3.80 ;
        RECT  19.85 3.15 20.75 5.00 ;
        RECT  20.20 3.10 20.70 9.60 ;
        RECT  20.00 3.15 20.70 9.60 ;
        RECT  20.20 3.10 20.75 5.95 ;
        RECT  20.00 3.15 20.75 5.95 ;
        RECT  20.20 3.10 20.90 3.80 ;
        RECT  19.85 3.15 20.90 3.80 ;
        RECT  20.20 3.10 22.10 3.65 ;
        RECT  21.40 2.45 22.10 3.65 ;
        RECT  7.90 3.15 22.10 3.65 ;
        RECT  20.00 5.45 23.35 5.95 ;
        RECT  22.85 5.45 23.35 9.60 ;
        RECT  22.85 7.10 23.55 9.60 ;
        RECT  22.85 8.90 23.75 9.60 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.57 ;
        PORT
        LAYER M1M ;
        RECT  22.65 4.10 23.55 5.00 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.57 ;
        PORT
        LAYER M1M ;
        RECT  18.45 4.10 19.35 5.00 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.57 ;
        PORT
        LAYER M1M ;
        RECT  14.20 4.10 15.15 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.57 ;
        PORT
        LAYER M1M ;
        RECT  17.05 4.10 17.95 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.35 3.95 6.30 ;
        RECT  3.05 5.60 4.25 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.35 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.40 1.15 11.00 ;
        RECT  1.85 10.40 2.55 11.00 ;
        RECT  4.20 7.70 4.90 11.00 ;
        RECT  2.80 7.70 6.30 8.40 ;
        RECT  7.95 7.70 8.65 11.00 ;
        RECT  6.55 10.40 10.05 11.00 ;
        RECT  10.30 7.70 12.40 8.40 ;
        RECT  11.70 7.70 12.40 11.00 ;
        RECT  0.00 11.00 26.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 2.00 1.20 4.80 ;
        RECT  2.05 2.00 2.75 4.50 ;
        RECT  9.50 2.00 13.50 2.65 ;
        RECT  17.85 2.00 18.55 2.70 ;
        RECT  22.90 2.00 26.15 3.65 ;
        RECT  24.00 2.00 26.15 3.80 ;
        RECT  0.00 0.00 26.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  12.15 6.40 18.00 6.70 ;
        RECT  1.80 6.75 2.30 9.75 ;
        RECT  1.80 9.05 3.55 9.75 ;
        RECT  6.80 6.75 7.30 9.75 ;
        RECT  5.55 9.05 7.30 9.75 ;
        RECT  9.30 6.75 9.80 9.75 ;
        RECT  9.30 9.05 11.05 9.75 ;
        RECT  12.15 6.20 12.65 7.25 ;
        RECT  1.80 6.75 12.65 7.25 ;
        RECT  13.25 7.15 13.95 10.55 ;
        RECT  14.60 6.20 15.10 9.25 ;
        RECT  12.15 6.20 15.10 6.70 ;
        RECT  14.60 6.40 15.30 9.25 ;
        RECT  15.95 7.35 16.65 10.55 ;
        RECT  14.60 6.40 18.00 6.90 ;
        RECT  17.30 6.40 18.00 9.60 ;
        RECT  18.65 6.40 19.35 10.55 ;
        RECT  21.35 6.40 22.05 10.55 ;
        RECT  24.60 7.15 25.30 10.55 ;
        RECT  13.25 10.05 25.30 10.55 ;
    END
END AN322X2
MACRO AN322X4
    CLASS CORE ;
    FOREIGN AN322X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 50.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  21.85 2.45 22.55 4.80 ;
        RECT  13.55 4.10 22.55 4.80 ;
        RECT  29.95 3.10 30.45 4.80 ;
        RECT  13.55 4.30 30.45 4.80 ;
        RECT  35.15 2.45 35.85 3.80 ;
        RECT  36.65 3.10 37.55 5.00 ;
        RECT  37.05 3.10 37.55 9.60 ;
        RECT  37.05 6.85 37.75 9.60 ;
        RECT  39.75 6.85 40.45 9.60 ;
        RECT  29.95 3.10 41.05 3.80 ;
        RECT  42.45 6.85 43.15 9.60 ;
        RECT  45.15 6.85 45.85 9.60 ;
        RECT  37.05 6.85 48.55 7.35 ;
        RECT  47.85 6.85 48.55 9.60 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 11.20 ;
        PORT
        LAYER M1M ;
        RECT  40.85 5.35 41.75 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 11.20 ;
        PORT
        LAYER M1M ;
        RECT  43.65 5.35 44.55 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 11.20 ;
        PORT
        LAYER M1M ;
        RECT  29.65 5.35 30.55 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 11.20 ;
        PORT
        LAYER M1M ;
        RECT  26.85 5.35 27.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.40 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.10 1.15 11.00 ;
        RECT  3.15 6.50 3.85 11.00 ;
        RECT  5.85 6.50 6.55 11.00 ;
        RECT  8.55 7.80 9.25 11.00 ;
        RECT  11.25 7.80 11.95 11.00 ;
        RECT  13.95 7.80 14.65 11.00 ;
        RECT  16.65 7.80 17.35 11.00 ;
        RECT  19.35 7.80 20.05 11.00 ;
        RECT  0.00 11.00 50.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 9.25 3.80 ;
        RECT  10.05 2.00 10.75 4.15 ;
        RECT  23.35 2.00 26.80 3.80 ;
        RECT  27.60 2.00 28.30 3.80 ;
        RECT  42.70 2.00 43.40 3.80 ;
        RECT  44.20 2.00 49.95 3.80 ;
        RECT  0.00 0.00 50.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 5.55 2.50 10.55 ;
        RECT  4.50 5.55 5.20 10.55 ;
        RECT  1.80 5.55 7.90 6.05 ;
        RECT  7.20 5.55 7.90 10.55 ;
        RECT  9.90 6.85 10.60 10.55 ;
        RECT  12.60 6.85 13.30 10.55 ;
        RECT  15.30 6.85 16.00 10.55 ;
        RECT  18.00 6.85 18.70 10.55 ;
        RECT  7.20 6.85 21.40 7.35 ;
        RECT  20.70 6.85 21.40 10.55 ;
        RECT  22.05 6.85 22.75 9.60 ;
        RECT  23.40 7.85 24.10 10.55 ;
        RECT  24.75 6.85 25.45 9.60 ;
        RECT  26.10 7.85 26.80 10.55 ;
        RECT  27.45 6.85 28.15 9.60 ;
        RECT  28.80 7.85 29.50 10.55 ;
        RECT  30.15 6.85 30.85 9.60 ;
        RECT  31.50 7.85 32.20 10.55 ;
        RECT  32.85 6.85 33.55 9.60 ;
        RECT  34.20 7.90 34.90 10.55 ;
        RECT  20.70 10.05 34.90 10.55 ;
        RECT  22.05 6.85 36.40 7.35 ;
        RECT  35.70 6.85 36.40 10.55 ;
        RECT  38.40 7.90 39.10 10.55 ;
        RECT  41.10 7.90 41.80 10.55 ;
        RECT  43.80 7.90 44.50 10.55 ;
        RECT  46.50 7.90 47.20 10.55 ;
        RECT  49.20 7.10 49.90 10.55 ;
        RECT  35.70 10.05 49.90 10.55 ;
    END
END AN322X4
MACRO AN32X1
    CLASS CORE ;
    FOREIGN AN32X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  3.80 2.45 4.50 4.85 ;
        RECT  3.80 4.35 6.55 4.85 ;
        RECT  6.05 4.35 6.55 9.60 ;
        RECT  5.85 7.20 6.55 9.60 ;
        RECT  5.85 8.00 6.75 8.90 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.35 5.35 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.35 3.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.35 2.60 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.20 1.15 11.00 ;
        RECT  3.15 8.05 3.85 11.00 ;
        RECT  0.00 11.00 8.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 4.20 ;
        RECT  6.30 2.00 7.00 3.85 ;
        RECT  0.00 0.00 8.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 7.05 2.50 10.55 ;
        RECT  1.80 7.05 5.20 7.55 ;
        RECT  4.50 7.05 5.20 10.55 ;
        RECT  7.20 7.20 7.90 10.55 ;
        RECT  4.50 10.05 7.90 10.55 ;
    END
END AN32X1
MACRO AN32X2
    CLASS CORE ;
    FOREIGN AN32X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  6.50 4.35 13.35 4.55 ;
        RECT  8.85 2.45 9.55 4.85 ;
        RECT  8.85 3.85 9.90 4.85 ;
        RECT  6.50 3.85 9.90 4.55 ;
        RECT  9.95 7.05 10.65 9.60 ;
        RECT  9.95 7.05 13.35 7.55 ;
        RECT  8.85 4.35 13.35 4.85 ;
        RECT  12.85 4.35 13.35 9.60 ;
        RECT  12.65 7.05 13.35 9.60 ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.20 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.35 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.20 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.20 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.40 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 8.05 2.55 11.00 ;
        RECT  4.55 8.05 5.25 11.00 ;
        RECT  7.25 8.05 7.95 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 2.20 4.70 ;
        RECT  3.00 2.00 3.70 4.50 ;
        RECT  11.70 2.00 12.40 3.85 ;
        RECT  13.20 2.00 14.95 3.80 ;
        RECT  13.80 2.00 14.95 4.70 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.50 7.05 1.20 10.55 ;
        RECT  3.20 7.05 3.90 10.55 ;
        RECT  5.90 7.05 6.60 10.55 ;
        RECT  0.50 7.05 9.30 7.55 ;
        RECT  8.60 7.05 9.30 10.55 ;
        RECT  11.30 8.05 12.00 10.55 ;
        RECT  14.00 7.15 14.70 10.55 ;
        RECT  8.60 10.05 14.70 10.55 ;
    END
END AN32X2
MACRO AN32X4
    CLASS CORE ;
    FOREIGN AN32X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 29.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.55 4.10 19.35 4.80 ;
        RECT  18.45 4.10 19.35 6.30 ;
        RECT  18.90 2.45 19.30 9.60 ;
        RECT  18.60 4.10 19.30 9.60 ;
        RECT  18.90 2.45 19.35 7.25 ;
        RECT  18.60 4.10 19.35 7.25 ;
        RECT  18.90 2.45 19.60 4.50 ;
        RECT  21.30 6.75 22.00 9.60 ;
        RECT  18.90 3.80 24.10 4.50 ;
        RECT  10.55 4.10 24.10 4.50 ;
        RECT  24.00 6.75 24.70 9.60 ;
        RECT  18.60 6.75 27.40 7.25 ;
        RECT  26.70 6.75 27.40 9.60 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 8.40 ;
        PORT
        LAYER M1M ;
        RECT  21.25 5.40 22.15 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 8.40 ;
        PORT
        LAYER M1M ;
        RECT  25.45 5.40 26.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.35 13.75 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.35 9.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.40 7.70 3.10 11.00 ;
        RECT  5.10 7.70 5.80 11.00 ;
        RECT  7.80 7.70 8.50 11.00 ;
        RECT  10.50 7.70 11.20 11.00 ;
        RECT  13.20 7.70 13.90 11.00 ;
        RECT  15.90 7.70 16.60 11.00 ;
        RECT  0.00 11.00 29.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 6.10 4.50 ;
        RECT  7.05 2.00 7.75 4.40 ;
        RECT  21.25 2.00 26.45 2.15 ;
        RECT  25.75 2.00 26.45 4.30 ;
        RECT  27.25 2.00 28.95 4.40 ;
        RECT  0.00 0.00 29.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.05 6.75 1.75 10.55 ;
        RECT  3.75 6.75 4.45 10.55 ;
        RECT  6.45 6.75 7.15 10.55 ;
        RECT  9.15 6.75 9.85 10.55 ;
        RECT  11.85 6.75 12.55 10.55 ;
        RECT  14.55 6.75 15.25 10.55 ;
        RECT  1.05 6.75 17.95 7.25 ;
        RECT  17.25 6.75 17.95 10.55 ;
        RECT  19.95 7.70 20.65 10.55 ;
        RECT  22.65 7.70 23.35 10.55 ;
        RECT  25.35 7.70 26.05 10.55 ;
        RECT  28.05 7.70 28.75 10.55 ;
        RECT  17.25 10.05 28.75 10.55 ;
    END
END AN32X4
MACRO AN331X1
    CLASS CORE ;
    FOREIGN AN331X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  5.80 2.45 6.30 3.65 ;
        RECT  3.80 2.45 6.30 3.15 ;
        RECT  10.25 6.70 10.95 10.20 ;
        RECT  10.50 2.90 11.20 3.65 ;
        RECT  5.80 3.15 11.90 3.65 ;
        RECT  11.40 3.15 11.90 7.60 ;
        RECT  10.25 6.70 12.35 7.60 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  10.05 4.10 10.95 5.00 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  5.85 4.10 6.75 5.00 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  7.25 4.10 8.15 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.55 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 3.95 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  1.65 4.10 2.55 5.00 ;
        RECT  1.85 4.10 2.55 5.55 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.80 8.20 1.50 11.00 ;
        RECT  3.50 6.95 4.20 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.70 ;
        RECT  9.00 2.00 9.70 2.70 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.15 6.00 2.85 10.55 ;
        RECT  2.15 6.00 5.55 6.50 ;
        RECT  4.85 6.00 5.55 10.55 ;
        RECT  6.20 6.00 6.90 9.60 ;
        RECT  7.55 6.95 8.25 10.55 ;
        RECT  4.85 10.05 8.25 10.55 ;
        RECT  6.20 6.00 9.60 6.50 ;
        RECT  8.90 6.00 9.60 10.55 ;
    END
END AN331X1
MACRO AN331X2
    CLASS CORE ;
    FOREIGN AN331X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 29.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  7.90 2.45 8.60 4.80 ;
        RECT  5.55 4.10 8.60 4.80 ;
        RECT  7.90 3.15 15.00 3.65 ;
        RECT  14.30 2.45 15.00 4.80 ;
        RECT  14.30 4.10 17.35 4.80 ;
        RECT  21.65 2.70 22.35 4.80 ;
        RECT  14.30 4.30 24.55 4.80 ;
        RECT  24.05 4.30 24.55 6.30 ;
        RECT  24.05 5.40 24.95 6.30 ;
        RECT  24.05 5.80 26.35 6.30 ;
        RECT  25.85 5.80 26.35 9.60 ;
        RECT  25.85 8.90 27.60 9.60 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  22.65 5.40 23.55 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  18.40 5.40 19.35 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.35 3.95 6.30 ;
        RECT  3.05 5.60 4.25 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.35 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.40 1.15 11.00 ;
        RECT  1.85 10.40 2.55 11.00 ;
        RECT  4.20 7.70 4.90 11.00 ;
        RECT  2.80 7.70 6.30 8.40 ;
        RECT  7.95 7.70 8.65 11.00 ;
        RECT  6.55 10.40 10.05 11.00 ;
        RECT  10.30 7.70 12.40 8.40 ;
        RECT  11.70 7.70 12.40 11.00 ;
        RECT  0.00 11.00 29.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 2.00 1.20 4.80 ;
        RECT  2.05 2.00 2.75 4.50 ;
        RECT  9.50 2.00 13.50 2.65 ;
        RECT  20.15 2.00 20.85 3.80 ;
        RECT  23.15 2.00 28.95 3.80 ;
        RECT  25.10 2.00 28.95 4.90 ;
        RECT  0.00 0.00 29.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 6.75 2.30 9.75 ;
        RECT  1.80 9.05 3.55 9.75 ;
        RECT  6.80 6.75 7.30 9.75 ;
        RECT  5.55 9.05 7.30 9.75 ;
        RECT  9.30 6.75 9.80 9.75 ;
        RECT  9.30 9.05 11.05 9.75 ;
        RECT  13.25 7.70 13.95 10.55 ;
        RECT  15.85 6.75 16.35 9.60 ;
        RECT  14.60 8.90 16.35 9.60 ;
        RECT  17.00 7.70 17.70 10.55 ;
        RECT  18.35 6.75 18.85 9.60 ;
        RECT  18.35 8.90 20.10 9.60 ;
        RECT  20.75 7.70 21.45 10.55 ;
        RECT  1.80 6.75 23.85 7.25 ;
        RECT  23.35 6.75 23.85 9.60 ;
        RECT  22.10 8.90 23.85 9.60 ;
        RECT  24.50 7.70 25.20 10.55 ;
        RECT  28.25 7.40 28.95 10.55 ;
        RECT  13.25 10.05 28.95 10.55 ;
    END
END AN331X2
MACRO AN331X4
    CLASS CORE ;
    FOREIGN AN331X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 50.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  21.85 2.45 22.55 4.85 ;
        RECT  13.55 4.10 22.55 4.85 ;
        RECT  42.10 2.45 42.80 4.85 ;
        RECT  33.80 4.10 42.80 4.85 ;
        RECT  42.30 6.85 43.00 9.60 ;
        RECT  13.55 4.35 44.15 4.85 ;
        RECT  43.65 4.35 44.15 7.35 ;
        RECT  43.65 5.40 44.55 7.35 ;
        RECT  45.00 6.85 45.70 9.60 ;
        RECT  42.30 6.85 48.40 7.35 ;
        RECT  47.70 6.85 48.40 10.55 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  42.25 5.40 43.15 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  35.25 5.40 36.15 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  31.00 5.40 31.95 6.40 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  28.25 5.40 29.15 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.40 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.10 1.15 11.00 ;
        RECT  3.15 6.50 3.85 11.00 ;
        RECT  5.85 6.50 6.55 11.00 ;
        RECT  8.55 7.80 9.25 11.00 ;
        RECT  11.25 7.80 11.95 11.00 ;
        RECT  13.95 7.80 14.65 11.00 ;
        RECT  16.65 7.80 17.35 11.00 ;
        RECT  19.35 7.80 20.05 11.00 ;
        RECT  49.25 9.55 49.95 11.00 ;
        RECT  0.00 11.00 50.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 9.25 3.80 ;
        RECT  10.05 2.00 10.75 4.15 ;
        RECT  23.35 2.00 29.50 3.80 ;
        RECT  30.30 2.00 31.00 3.90 ;
        RECT  43.45 2.00 44.15 3.90 ;
        RECT  44.95 2.00 49.95 4.75 ;
        RECT  0.00 0.00 50.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 5.55 2.50 10.55 ;
        RECT  4.50 5.55 5.20 10.55 ;
        RECT  1.80 5.55 7.90 6.05 ;
        RECT  7.20 5.55 7.90 10.55 ;
        RECT  9.90 6.85 10.60 10.55 ;
        RECT  12.60 6.85 13.30 10.55 ;
        RECT  15.30 6.85 16.00 10.55 ;
        RECT  18.00 6.85 18.70 10.55 ;
        RECT  7.20 6.85 21.40 7.35 ;
        RECT  20.70 6.85 21.40 10.55 ;
        RECT  22.05 6.85 22.75 9.60 ;
        RECT  23.40 7.85 24.10 10.55 ;
        RECT  24.75 6.85 25.45 9.60 ;
        RECT  26.10 7.85 26.80 10.55 ;
        RECT  27.45 6.85 28.15 9.60 ;
        RECT  28.80 7.85 29.50 10.55 ;
        RECT  30.15 6.85 30.85 9.60 ;
        RECT  31.50 7.85 32.20 10.55 ;
        RECT  32.85 6.85 33.55 9.60 ;
        RECT  34.20 7.90 34.90 10.55 ;
        RECT  35.55 6.85 36.25 9.60 ;
        RECT  36.90 7.90 37.60 10.55 ;
        RECT  38.25 6.85 38.95 9.60 ;
        RECT  39.60 7.90 40.30 10.55 ;
        RECT  20.70 10.05 40.30 10.55 ;
        RECT  22.05 6.85 41.65 7.35 ;
        RECT  40.95 6.85 41.65 10.55 ;
        RECT  43.65 7.90 44.35 10.55 ;
        RECT  46.35 7.90 47.05 10.55 ;
        RECT  40.95 10.05 47.05 10.55 ;
    END
END AN331X4
MACRO AN332X1
    CLASS CORE ;
    FOREIGN AN332X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  3.80 3.15 13.75 3.50 ;
        RECT  6.30 2.80 6.80 3.65 ;
        RECT  3.80 2.80 6.80 3.50 ;
        RECT  10.45 5.45 10.95 9.60 ;
        RECT  10.25 6.40 10.95 9.60 ;
        RECT  12.00 2.60 12.70 3.65 ;
        RECT  12.00 2.80 13.75 3.65 ;
        RECT  6.30 3.15 13.75 3.65 ;
        RECT  12.80 2.80 13.30 5.95 ;
        RECT  10.45 5.45 13.30 5.95 ;
        RECT  12.80 2.80 13.75 3.70 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  11.45 4.10 12.35 5.00 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  10.05 4.10 10.95 5.00 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  5.85 4.10 6.75 5.00 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  7.20 4.10 7.90 5.65 ;
        RECT  7.20 4.10 8.15 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.55 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 3.95 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  1.65 4.10 2.55 5.00 ;
        RECT  1.85 4.10 2.55 5.65 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.80 8.20 1.50 11.00 ;
        RECT  3.50 7.05 4.20 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.80 ;
        RECT  9.50 2.00 10.20 2.70 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.15 6.10 2.85 10.55 ;
        RECT  2.15 6.10 5.55 6.60 ;
        RECT  4.85 6.10 5.55 10.55 ;
        RECT  6.20 6.10 6.90 9.60 ;
        RECT  7.55 7.05 8.25 10.55 ;
        RECT  4.85 10.05 8.25 10.55 ;
        RECT  6.20 6.10 9.60 6.60 ;
        RECT  8.90 6.10 9.60 10.55 ;
        RECT  11.60 6.85 12.30 10.55 ;
        RECT  8.90 10.05 12.30 10.55 ;
    END
END AN332X1
MACRO AN332X2
    CLASS CORE ;
    FOREIGN AN332X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 33.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  7.90 2.45 8.60 4.80 ;
        RECT  5.55 4.10 8.60 4.80 ;
        RECT  14.30 2.45 15.00 4.80 ;
        RECT  14.30 4.10 17.35 4.80 ;
        RECT  25.45 5.40 26.35 6.30 ;
        RECT  25.85 4.30 26.35 9.60 ;
        RECT  25.85 8.90 27.60 9.60 ;
        RECT  25.85 6.75 30.10 7.25 ;
        RECT  29.60 6.75 30.10 9.60 ;
        RECT  29.60 8.90 31.35 9.60 ;
        RECT  31.95 3.80 32.70 4.80 ;
        RECT  32.20 2.45 32.70 4.80 ;
        RECT  5.55 4.30 32.70 4.80 ;
        RECT  32.20 2.45 33.15 3.15 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.60 ;
        PORT
        LAYER M1M ;
        RECT  31.05 5.40 32.20 6.30 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.60 ;
        PORT
        LAYER M1M ;
        RECT  26.85 5.40 27.75 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  18.40 5.40 19.35 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.35 3.95 6.30 ;
        RECT  3.05 5.60 4.25 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.35 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.40 1.15 11.00 ;
        RECT  1.85 10.40 2.55 11.00 ;
        RECT  4.20 7.70 4.90 11.00 ;
        RECT  2.80 7.70 6.30 8.40 ;
        RECT  7.95 7.70 8.65 11.00 ;
        RECT  6.55 10.40 10.05 11.00 ;
        RECT  10.30 7.70 12.40 8.40 ;
        RECT  11.70 7.70 12.40 11.00 ;
        RECT  0.00 11.00 33.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 2.00 1.20 4.80 ;
        RECT  2.05 2.00 2.75 4.50 ;
        RECT  9.50 2.00 13.50 3.80 ;
        RECT  20.15 2.00 20.85 3.80 ;
        RECT  21.65 2.00 28.80 3.80 ;
        RECT  29.60 2.00 30.30 3.85 ;
        RECT  0.00 0.00 33.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 6.75 2.30 9.75 ;
        RECT  1.80 9.05 3.55 9.75 ;
        RECT  6.80 6.75 7.30 9.75 ;
        RECT  5.55 9.05 7.30 9.75 ;
        RECT  9.30 6.75 9.80 9.75 ;
        RECT  9.30 9.05 11.05 9.75 ;
        RECT  13.25 7.70 13.95 10.55 ;
        RECT  15.85 6.75 16.35 9.60 ;
        RECT  14.60 8.90 16.35 9.60 ;
        RECT  17.00 7.70 17.70 10.55 ;
        RECT  18.35 6.75 18.85 9.60 ;
        RECT  18.35 8.90 20.10 9.60 ;
        RECT  20.75 7.70 21.45 10.55 ;
        RECT  1.80 6.75 23.85 7.25 ;
        RECT  23.35 6.75 23.85 9.60 ;
        RECT  22.10 8.90 23.85 9.60 ;
        RECT  24.50 7.70 25.20 10.55 ;
        RECT  28.25 7.70 28.95 10.55 ;
        RECT  30.60 7.40 32.70 8.10 ;
        RECT  32.00 7.40 32.70 10.55 ;
        RECT  13.25 10.05 32.70 10.55 ;
    END
END AN332X2
MACRO AN332X4
    CLASS CORE ;
    FOREIGN AN332X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 56.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  42.25 5.40 43.15 6.30 ;
        RECT  21.85 2.45 22.55 4.85 ;
        RECT  13.55 4.10 22.55 4.85 ;
        RECT  33.80 4.10 42.80 4.85 ;
        RECT  42.10 2.45 42.80 4.85 ;
        RECT  13.55 4.35 42.80 4.85 ;
        RECT  42.30 2.45 42.80 9.60 ;
        RECT  42.25 2.45 42.80 6.30 ;
        RECT  42.30 5.40 43.00 9.60 ;
        RECT  42.30 5.40 43.15 7.35 ;
        RECT  45.00 6.85 45.70 9.60 ;
        RECT  42.10 3.10 48.00 3.80 ;
        RECT  47.70 6.85 48.40 9.60 ;
        RECT  50.40 6.85 51.10 9.60 ;
        RECT  42.30 6.85 53.80 7.35 ;
        RECT  53.10 6.85 53.80 9.60 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 11.20 ;
        PORT
        LAYER M1M ;
        RECT  46.45 5.35 47.35 6.30 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 11.20 ;
        PORT
        LAYER M1M ;
        RECT  49.25 4.10 50.15 5.00 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  33.85 5.40 34.75 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  31.00 5.40 31.95 6.40 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  28.25 5.40 29.15 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.40 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.10 1.15 11.00 ;
        RECT  3.15 6.50 3.85 11.00 ;
        RECT  5.85 6.50 6.55 11.00 ;
        RECT  8.55 7.80 9.25 11.00 ;
        RECT  11.25 7.80 11.95 11.00 ;
        RECT  13.95 7.80 14.65 11.00 ;
        RECT  16.65 7.80 17.35 11.00 ;
        RECT  19.35 7.80 20.05 11.00 ;
        RECT  0.00 11.00 56.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 9.25 3.80 ;
        RECT  10.05 2.00 10.75 4.15 ;
        RECT  23.35 2.00 29.50 3.80 ;
        RECT  30.30 2.00 31.00 3.90 ;
        RECT  49.65 2.00 50.35 3.65 ;
        RECT  51.20 2.00 55.50 3.85 ;
        RECT  0.00 0.00 56.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 5.55 2.50 10.55 ;
        RECT  4.50 5.55 5.20 10.55 ;
        RECT  1.80 5.55 7.90 6.05 ;
        RECT  7.20 5.55 7.90 10.55 ;
        RECT  9.90 6.85 10.60 10.55 ;
        RECT  12.60 6.85 13.30 10.55 ;
        RECT  15.30 6.85 16.00 10.55 ;
        RECT  18.00 6.85 18.70 10.55 ;
        RECT  7.20 6.85 21.40 7.35 ;
        RECT  20.70 6.85 21.40 10.55 ;
        RECT  22.05 6.85 22.75 9.60 ;
        RECT  23.40 7.85 24.10 10.55 ;
        RECT  24.75 6.85 25.45 9.60 ;
        RECT  26.10 7.85 26.80 10.55 ;
        RECT  27.45 6.85 28.15 9.60 ;
        RECT  28.80 7.85 29.50 10.55 ;
        RECT  30.15 6.85 30.85 9.60 ;
        RECT  31.50 7.85 32.20 10.55 ;
        RECT  32.85 6.85 33.55 9.60 ;
        RECT  34.20 7.90 34.90 10.55 ;
        RECT  35.55 6.85 36.25 9.60 ;
        RECT  36.90 7.90 37.60 10.55 ;
        RECT  38.25 6.85 38.95 9.60 ;
        RECT  39.60 7.90 40.30 10.55 ;
        RECT  20.70 10.05 40.30 10.55 ;
        RECT  22.05 6.85 41.65 7.35 ;
        RECT  40.95 6.85 41.65 10.55 ;
        RECT  43.65 7.90 44.35 10.55 ;
        RECT  46.35 7.90 47.05 10.55 ;
        RECT  49.05 7.90 49.75 10.55 ;
        RECT  51.75 7.90 52.45 10.55 ;
        RECT  54.45 7.10 55.15 10.55 ;
        RECT  40.95 10.05 55.15 10.55 ;
    END
END AN332X4
MACRO AN333X1
    CLASS CORE ;
    FOREIGN AN333X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  3.80 3.15 15.15 3.50 ;
        RECT  6.30 2.80 6.80 3.65 ;
        RECT  3.80 2.80 6.80 3.50 ;
        RECT  10.25 5.45 10.95 9.60 ;
        RECT  12.95 5.45 13.65 10.20 ;
        RECT  13.10 2.80 15.15 3.65 ;
        RECT  6.30 3.15 15.15 3.65 ;
        RECT  14.20 2.80 14.70 5.95 ;
        RECT  10.25 5.45 14.70 5.95 ;
        RECT  14.20 2.80 15.15 3.70 ;
        END
    END Q
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  10.05 4.10 10.95 5.00 ;
        END
    END J
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  11.40 4.10 12.35 5.00 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  12.85 4.10 13.75 5.00 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  5.85 4.10 6.75 5.00 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  7.20 4.10 7.90 5.65 ;
        RECT  7.20 4.10 8.15 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.55 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 3.95 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  1.65 4.10 2.55 5.00 ;
        RECT  1.85 4.10 2.55 5.65 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.80 8.20 1.50 11.00 ;
        RECT  3.50 7.05 4.20 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.80 ;
        RECT  9.60 2.00 10.30 2.70 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.15 6.10 2.85 10.55 ;
        RECT  2.15 6.10 5.55 6.60 ;
        RECT  4.85 6.10 5.55 10.55 ;
        RECT  6.20 6.10 6.90 9.60 ;
        RECT  7.55 7.05 8.25 10.55 ;
        RECT  4.85 10.05 8.25 10.55 ;
        RECT  6.20 6.10 9.60 6.60 ;
        RECT  8.90 6.10 9.60 10.55 ;
        RECT  11.60 6.40 12.30 10.55 ;
        RECT  8.90 10.05 12.30 10.55 ;
    END
END AN333X1
MACRO AN333X2
    CLASS CORE ;
    FOREIGN AN333X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 37.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  7.90 2.45 8.60 4.80 ;
        RECT  5.55 4.10 8.60 4.80 ;
        RECT  14.30 2.45 15.00 4.80 ;
        RECT  14.30 4.10 17.35 4.80 ;
        RECT  25.85 6.75 26.35 9.60 ;
        RECT  25.85 8.90 27.60 9.60 ;
        RECT  28.25 5.40 29.15 6.30 ;
        RECT  28.65 4.30 29.15 7.25 ;
        RECT  29.60 6.75 30.10 9.60 ;
        RECT  29.60 8.90 31.35 9.60 ;
        RECT  25.85 6.75 33.85 7.25 ;
        RECT  33.35 6.75 33.85 9.60 ;
        RECT  31.70 4.10 34.75 4.80 ;
        RECT  34.05 2.45 34.75 4.80 ;
        RECT  5.55 4.30 34.75 4.80 ;
        RECT  33.35 8.90 35.10 9.60 ;
        END
    END Q
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  26.85 5.40 27.75 6.30 ;
        END
    END J
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  29.65 5.40 30.55 6.30 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  33.85 5.40 34.75 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  18.40 5.40 19.35 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.35 3.95 6.30 ;
        RECT  3.05 5.60 4.25 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.35 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.40 1.15 11.00 ;
        RECT  1.85 10.40 2.55 11.00 ;
        RECT  4.20 7.70 4.90 11.00 ;
        RECT  2.80 7.70 6.30 8.40 ;
        RECT  7.95 7.70 8.65 11.00 ;
        RECT  6.55 10.40 10.05 11.00 ;
        RECT  10.30 7.70 12.40 8.40 ;
        RECT  11.70 7.70 12.40 11.00 ;
        RECT  0.00 11.00 37.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 2.00 1.20 4.80 ;
        RECT  2.05 2.00 2.75 4.50 ;
        RECT  9.50 2.00 13.50 3.80 ;
        RECT  20.15 2.00 20.85 3.80 ;
        RECT  21.65 2.00 27.40 3.80 ;
        RECT  28.20 2.00 28.90 3.85 ;
        RECT  35.55 2.00 37.35 4.70 ;
        RECT  0.00 0.00 37.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 6.75 2.30 9.75 ;
        RECT  1.80 9.05 3.55 9.75 ;
        RECT  6.80 6.75 7.30 9.75 ;
        RECT  5.55 9.05 7.30 9.75 ;
        RECT  9.30 6.75 9.80 9.75 ;
        RECT  9.30 9.05 11.05 9.75 ;
        RECT  13.25 7.70 13.95 10.55 ;
        RECT  15.85 6.75 16.35 9.60 ;
        RECT  14.60 8.90 16.35 9.60 ;
        RECT  17.00 7.70 17.70 10.55 ;
        RECT  18.35 6.75 18.85 9.60 ;
        RECT  18.35 8.90 20.10 9.60 ;
        RECT  20.75 7.70 21.45 10.55 ;
        RECT  1.80 6.75 23.85 7.25 ;
        RECT  23.35 6.75 23.85 9.60 ;
        RECT  22.10 8.90 23.85 9.60 ;
        RECT  24.50 7.70 25.20 10.55 ;
        RECT  28.25 7.70 28.95 10.55 ;
        RECT  32.00 7.70 32.70 10.55 ;
        RECT  35.75 7.40 36.45 10.55 ;
        RECT  13.25 10.05 36.45 10.55 ;
    END
END AN333X2
MACRO AN333X4
    CLASS CORE ;
    FOREIGN AN333X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 63.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  42.25 5.40 43.15 6.30 ;
        RECT  21.85 2.45 22.55 4.85 ;
        RECT  13.55 4.10 22.55 4.85 ;
        RECT  42.10 2.45 42.80 4.85 ;
        RECT  42.30 2.45 42.80 9.60 ;
        RECT  42.25 2.45 42.80 6.30 ;
        RECT  42.30 5.40 43.00 9.60 ;
        RECT  42.30 5.40 43.15 7.35 ;
        RECT  45.00 6.85 45.70 9.60 ;
        RECT  47.70 6.85 48.40 9.60 ;
        RECT  33.80 4.10 51.10 4.85 ;
        RECT  13.55 4.35 51.10 4.85 ;
        RECT  50.40 6.85 51.10 9.60 ;
        RECT  53.10 6.85 53.80 9.60 ;
        RECT  55.80 6.85 56.50 9.60 ;
        RECT  58.50 6.85 59.20 9.60 ;
        RECT  42.30 6.85 61.90 7.35 ;
        RECT  61.20 6.85 61.90 10.55 ;
        END
    END Q
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  54.85 5.40 55.75 6.30 ;
        END
    END J
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  52.05 5.35 52.95 6.30 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  49.25 5.40 50.15 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  33.85 5.40 34.75 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  31.00 5.40 31.95 6.40 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  28.25 5.40 29.15 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.40 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.10 1.15 11.00 ;
        RECT  3.15 6.50 3.85 11.00 ;
        RECT  5.85 6.50 6.55 11.00 ;
        RECT  8.55 7.80 9.25 11.00 ;
        RECT  11.25 7.80 11.95 11.00 ;
        RECT  13.95 7.80 14.65 11.00 ;
        RECT  16.65 7.80 17.35 11.00 ;
        RECT  19.35 7.80 20.05 11.00 ;
        RECT  0.00 11.00 63.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 9.25 3.80 ;
        RECT  10.05 2.00 10.75 4.15 ;
        RECT  23.35 2.00 29.50 3.80 ;
        RECT  30.30 2.00 31.00 3.90 ;
        RECT  53.90 2.00 54.60 3.90 ;
        RECT  55.45 2.00 62.50 3.85 ;
        RECT  0.00 0.00 63.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 5.55 2.50 10.55 ;
        RECT  4.50 5.55 5.20 10.55 ;
        RECT  1.80 5.55 7.90 6.05 ;
        RECT  7.20 5.55 7.90 10.55 ;
        RECT  9.90 6.85 10.60 10.55 ;
        RECT  12.60 6.85 13.30 10.55 ;
        RECT  15.30 6.85 16.00 10.55 ;
        RECT  18.00 6.85 18.70 10.55 ;
        RECT  7.20 6.85 21.40 7.35 ;
        RECT  20.70 6.85 21.40 10.55 ;
        RECT  22.05 6.85 22.75 9.60 ;
        RECT  23.40 7.85 24.10 10.55 ;
        RECT  24.75 6.85 25.45 9.60 ;
        RECT  26.10 7.85 26.80 10.55 ;
        RECT  27.45 6.85 28.15 9.60 ;
        RECT  28.80 7.85 29.50 10.55 ;
        RECT  30.15 6.85 30.85 9.60 ;
        RECT  31.50 7.85 32.20 10.55 ;
        RECT  32.85 6.85 33.55 9.60 ;
        RECT  34.20 7.90 34.90 10.55 ;
        RECT  35.55 6.85 36.25 9.60 ;
        RECT  36.90 7.90 37.60 10.55 ;
        RECT  38.25 6.85 38.95 9.60 ;
        RECT  39.60 7.90 40.30 10.55 ;
        RECT  20.70 10.05 40.30 10.55 ;
        RECT  22.05 6.85 41.65 7.35 ;
        RECT  40.95 6.85 41.65 10.55 ;
        RECT  43.65 7.90 44.35 10.55 ;
        RECT  46.35 7.90 47.05 10.55 ;
        RECT  49.05 7.90 49.75 10.55 ;
        RECT  51.75 7.90 52.45 10.55 ;
        RECT  54.45 7.90 55.15 10.55 ;
        RECT  57.15 7.90 57.85 10.55 ;
        RECT  59.85 7.90 60.55 10.55 ;
        RECT  40.95 10.05 60.55 10.55 ;
    END
END AN333X4
MACRO AN33X1
    CLASS CORE ;
    FOREIGN AN33X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  3.80 2.45 4.50 4.60 ;
        RECT  5.85 6.75 6.55 9.60 ;
        RECT  3.80 4.10 8.15 4.60 ;
        RECT  7.25 4.10 7.75 7.35 ;
        RECT  7.25 4.10 8.15 5.00 ;
        RECT  5.85 6.75 9.25 7.35 ;
        RECT  8.55 6.75 9.25 10.55 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.35 5.35 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.35 6.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.40 9.55 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.35 3.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.35 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.20 1.15 11.00 ;
        RECT  3.15 7.70 3.85 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 4.20 ;
        RECT  7.15 2.00 7.85 3.65 ;
        RECT  8.65 2.00 9.35 4.75 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 6.75 2.50 10.55 ;
        RECT  1.80 6.75 5.20 7.25 ;
        RECT  4.50 6.75 5.20 10.55 ;
        RECT  7.20 7.80 7.90 10.55 ;
        RECT  4.50 10.05 7.90 10.55 ;
    END
END AN33X1
MACRO AN33X2
    CLASS CORE ;
    FOREIGN AN33X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.00 2.45 8.70 4.55 ;
        RECT  10.05 3.85 10.55 9.60 ;
        RECT  10.05 6.85 10.65 9.60 ;
        RECT  9.95 7.45 10.65 9.60 ;
        RECT  5.75 3.85 10.95 4.55 ;
        RECT  10.05 5.40 10.95 6.30 ;
        RECT  12.65 6.85 13.35 9.60 ;
        RECT  10.05 6.85 16.05 7.35 ;
        RECT  15.35 6.85 16.05 9.60 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.35 9.55 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.65 6.40 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.35 15.15 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.35 8.15 6.35 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  4.00 5.35 5.35 6.35 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 7.75 2.55 11.00 ;
        RECT  4.55 7.75 5.25 11.00 ;
        RECT  7.25 7.75 7.95 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.55 2.00 1.25 4.75 ;
        RECT  2.15 2.00 2.85 4.30 ;
        RECT  13.85 2.00 14.55 4.30 ;
        RECT  15.35 2.00 17.75 4.75 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.50 6.80 1.20 10.55 ;
        RECT  3.20 6.80 3.90 10.55 ;
        RECT  5.90 6.80 6.60 10.55 ;
        RECT  0.50 6.80 9.30 7.30 ;
        RECT  8.60 6.80 9.30 10.55 ;
        RECT  11.30 7.80 12.00 10.55 ;
        RECT  14.00 7.80 14.70 10.55 ;
        RECT  16.70 7.80 17.40 10.55 ;
        RECT  8.60 10.05 17.40 10.55 ;
    END
END AN33X2
MACRO AN33X4
    CLASS CORE ;
    FOREIGN AN33X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 35.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  17.15 2.45 17.85 4.80 ;
        RECT  18.45 4.10 19.35 6.30 ;
        RECT  18.60 4.10 19.30 9.60 ;
        RECT  18.60 4.10 19.35 7.25 ;
        RECT  21.30 6.75 22.00 9.60 ;
        RECT  24.00 6.75 24.70 9.60 ;
        RECT  8.80 4.10 26.20 4.80 ;
        RECT  26.70 6.75 27.40 9.60 ;
        RECT  29.40 6.75 30.10 9.60 ;
        RECT  18.60 6.75 32.80 7.25 ;
        RECT  32.10 6.75 32.80 9.60 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  21.25 5.40 22.15 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  26.85 5.40 28.05 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  29.65 5.40 30.55 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.35 13.75 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  6.90 5.35 8.15 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.40 7.70 3.10 11.00 ;
        RECT  5.10 7.70 5.80 11.00 ;
        RECT  7.80 7.70 8.50 11.00 ;
        RECT  10.50 7.70 11.20 11.00 ;
        RECT  13.20 7.70 13.90 11.00 ;
        RECT  15.90 7.70 16.60 11.00 ;
        RECT  0.00 11.00 35.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 4.35 4.50 ;
        RECT  5.30 2.00 6.00 4.40 ;
        RECT  29.00 2.00 29.70 4.40 ;
        RECT  30.65 2.00 34.55 4.40 ;
        RECT  0.00 0.00 35.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.05 6.75 1.75 10.55 ;
        RECT  3.75 6.75 4.45 10.55 ;
        RECT  6.45 6.75 7.15 10.55 ;
        RECT  9.15 6.75 9.85 10.55 ;
        RECT  11.85 6.75 12.55 10.55 ;
        RECT  14.55 6.75 15.25 10.55 ;
        RECT  1.05 6.75 17.95 7.25 ;
        RECT  17.25 6.75 17.95 10.55 ;
        RECT  19.95 7.70 20.65 10.55 ;
        RECT  22.65 7.70 23.35 10.55 ;
        RECT  25.35 7.70 26.05 10.55 ;
        RECT  28.05 7.70 28.75 10.55 ;
        RECT  30.75 7.70 31.45 10.55 ;
        RECT  33.45 7.70 34.15 10.55 ;
        RECT  17.25 10.05 34.15 10.55 ;
    END
END AN33X4
MACRO AND2X1
    CLASS CORE ;
    FOREIGN AND2X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.15 3.15 4.85 3.85 ;
        RECT  4.35 3.15 4.85 9.40 ;
        RECT  4.15 7.70 4.85 9.40 ;
        RECT  4.15 8.00 5.35 8.90 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.10 9.90 1.80 11.00 ;
        RECT  2.80 7.70 3.50 11.00 ;
        RECT  0.00 11.00 5.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 2.00 3.50 3.85 ;
        RECT  0.00 0.00 5.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.15 1.15 4.95 ;
        RECT  1.10 6.75 1.80 9.25 ;
        RECT  0.45 4.45 3.90 4.95 ;
        RECT  3.00 4.45 3.50 7.25 ;
        RECT  1.10 6.75 3.50 7.25 ;
        RECT  3.00 4.45 3.90 5.15 ;
    END
END AND2X1
MACRO AND2X2
    CLASS CORE ;
    FOREIGN AND2X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.30 2.45 5.00 4.05 ;
        RECT  4.45 2.45 4.90 10.55 ;
        RECT  4.20 7.15 4.90 10.55 ;
        RECT  4.45 2.45 5.00 8.90 ;
        RECT  4.20 7.15 5.00 8.90 ;
        RECT  4.20 8.00 5.35 8.90 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.15 9.35 1.85 11.00 ;
        RECT  2.85 7.70 3.55 11.00 ;
        RECT  0.00 11.00 5.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.95 2.00 3.65 4.00 ;
        RECT  0.00 0.00 5.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.35 1.15 4.95 ;
        RECT  1.15 6.75 1.85 8.70 ;
        RECT  0.45 4.45 4.00 4.95 ;
        RECT  3.00 4.45 3.50 7.25 ;
        RECT  1.15 6.75 3.50 7.25 ;
        RECT  3.00 4.45 4.00 5.15 ;
    END
END AND2X2
MACRO AND2X3
    CLASS CORE ;
    FOREIGN AND2X3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.30 2.45 5.00 4.05 ;
        RECT  4.45 2.45 5.00 10.55 ;
        RECT  4.45 7.15 5.15 10.55 ;
        RECT  4.05 9.85 5.15 10.55 ;
        RECT  4.45 8.00 5.35 8.90 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 9.35 1.65 11.00 ;
        RECT  2.55 7.70 3.35 11.00 ;
        RECT  0.00 11.00 5.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.95 2.00 3.65 4.00 ;
        RECT  0.00 0.00 5.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.35 1.15 4.95 ;
        RECT  0.95 6.75 1.65 8.70 ;
        RECT  0.45 4.45 4.00 4.95 ;
        RECT  3.00 4.45 3.50 7.25 ;
        RECT  0.95 6.75 3.50 7.25 ;
        RECT  3.00 4.45 4.00 5.15 ;
    END
END AND2X3
MACRO AND2X4
    CLASS CORE ;
    FOREIGN AND2X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.30 2.45 5.00 4.05 ;
        RECT  4.45 2.45 4.95 10.55 ;
        RECT  4.20 7.15 4.95 10.55 ;
        RECT  4.45 2.45 5.00 6.30 ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.15 9.35 1.85 11.00 ;
        RECT  2.85 7.70 3.55 11.00 ;
        RECT  5.55 7.70 6.25 11.00 ;
        RECT  0.00 11.00 7.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.95 2.00 3.65 4.00 ;
        RECT  5.65 2.00 6.35 4.00 ;
        RECT  0.00 0.00 7.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.35 1.15 4.95 ;
        RECT  1.15 6.75 1.85 8.70 ;
        RECT  0.45 4.45 4.00 4.95 ;
        RECT  3.00 4.45 3.50 7.25 ;
        RECT  1.15 6.75 3.50 7.25 ;
        RECT  3.00 4.45 4.00 5.15 ;
    END
END AND2X4
MACRO AND3X1
    CLASS CORE ;
    FOREIGN AND3X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  5.35 3.55 6.35 4.25 ;
        RECT  5.85 3.55 6.35 9.30 ;
        RECT  5.85 6.70 6.75 9.30 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.70 2.50 11.00 ;
        RECT  0.45 10.10 2.95 11.00 ;
        RECT  4.35 7.70 5.20 11.00 ;
        RECT  0.00 11.00 7.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.80 2.00 4.50 4.00 ;
        RECT  0.00 0.00 7.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.40 1.15 4.95 ;
        RECT  0.45 6.75 1.15 8.50 ;
        RECT  3.15 6.75 3.85 8.50 ;
        RECT  0.45 4.45 4.90 4.95 ;
        RECT  4.40 4.45 4.90 7.25 ;
        RECT  0.45 6.75 4.90 7.25 ;
        RECT  4.40 5.50 5.40 6.20 ;
    END
END AND3X1
MACRO AND3X2
    CLASS CORE ;
    FOREIGN AND3X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  5.35 2.45 6.05 5.00 ;
        RECT  6.05 4.10 6.55 10.55 ;
        RECT  5.85 7.10 6.55 10.55 ;
        RECT  5.35 4.10 6.75 5.00 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.70 2.50 11.00 ;
        RECT  0.45 10.10 2.95 11.00 ;
        RECT  4.50 7.70 5.20 11.00 ;
        RECT  0.00 11.00 7.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.95 2.00 4.65 4.00 ;
        RECT  0.00 0.00 7.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.40 1.15 4.95 ;
        RECT  0.45 6.75 1.15 8.50 ;
        RECT  3.15 6.75 3.85 8.50 ;
        RECT  0.45 4.45 4.90 4.95 ;
        RECT  4.40 4.45 4.90 7.25 ;
        RECT  0.45 6.75 4.90 7.25 ;
        RECT  4.40 5.50 5.60 6.20 ;
    END
END AND3X2
MACRO AND3X3
    CLASS CORE ;
    FOREIGN AND3X3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  5.35 2.45 6.05 5.00 ;
        RECT  6.05 4.10 6.55 10.55 ;
        RECT  5.85 7.10 6.55 10.55 ;
        RECT  5.35 4.10 6.75 5.00 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.70 2.50 11.00 ;
        RECT  0.45 10.10 2.95 11.00 ;
        RECT  4.50 7.70 4.65 11.00 ;
        RECT  3.95 8.95 4.65 11.00 ;
        RECT  4.50 7.70 5.20 9.65 ;
        RECT  3.95 8.95 5.20 9.65 ;
        RECT  0.00 11.00 7.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.95 2.00 4.65 4.00 ;
        RECT  0.00 0.00 7.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.40 1.15 4.95 ;
        RECT  0.45 6.75 1.15 8.50 ;
        RECT  3.15 6.75 3.85 8.50 ;
        RECT  0.45 4.45 4.90 4.95 ;
        RECT  4.40 4.45 4.90 7.25 ;
        RECT  0.45 6.75 4.90 7.25 ;
        RECT  4.40 5.50 5.60 6.20 ;
    END
END AND3X3
MACRO AND3X4
    CLASS CORE ;
    FOREIGN AND3X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  6.05 2.45 6.15 10.55 ;
        RECT  5.35 2.45 6.15 5.00 ;
        RECT  6.05 4.10 6.55 10.55 ;
        RECT  5.85 7.10 6.55 10.55 ;
        RECT  5.35 4.10 6.75 5.00 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.70 2.50 11.00 ;
        RECT  0.45 10.10 2.50 11.00 ;
        RECT  2.95 9.20 3.65 11.00 ;
        RECT  4.50 7.70 5.20 9.90 ;
        RECT  2.95 9.20 5.20 9.90 ;
        RECT  0.00 11.00 7.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.95 2.00 4.65 4.00 ;
        RECT  0.00 0.00 7.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.30 1.15 4.95 ;
        RECT  0.45 6.75 1.15 8.40 ;
        RECT  3.15 6.75 3.85 8.40 ;
        RECT  0.45 4.45 4.90 4.95 ;
        RECT  4.40 4.45 4.90 7.25 ;
        RECT  0.45 6.75 4.90 7.25 ;
        RECT  4.40 5.50 5.60 6.20 ;
    END
END AND3X4
#MACRO AND4X1
#    CLASS CORE ;
#    FOREIGN AND4X1 0.00 0.00  ;
#    ORIGIN 0.00 0.00 ;
#    SIZE 11.20 BY 13.00 ;
#    SYMMETRY x y r90 ;
#    SITE core ;
#    PIN Q
#        DIRECTION OUTPUT ;
#        ANTENNADIFFAREA 1.0 ;
#        PORT
#        LAYER M1M ;
#        RECT  4.85 2.95 5.55 3.65 ;
#        RECT  5.05 2.95 5.55 5.90 ;
#        RECT  5.05 5.40 6.75 5.90 ;
#        RECT  5.65 5.40 6.35 10.55 ;
#        RECT  5.65 5.40 6.75 6.30 ;
#        END
#    END Q
#    PIN D
#        DIRECTION INPUT ;
#        ANTENNAGATEAREA 0.70 ;
#        PORT
#        LAYER M1M ;
#        RECT  8.65 5.40 9.55 6.30 ;
#        END
#    END D
#    PIN C
#        DIRECTION INPUT ;
#        ANTENNAGATEAREA 0.70 ;
#        PORT
#        LAYER M1M ;
#        RECT  10.05 4.10 10.95 5.00 ;
#        END
#    END C
#    PIN B
#        DIRECTION INPUT ;
#        ANTENNAGATEAREA 0.70 ;
#        PORT
#        LAYER M1M ;
#        RECT  1.65 4.10 2.55 5.00 ;
#        END
#    END B
#    PIN A
#        DIRECTION INPUT ;
#        ANTENNAGATEAREA 0.70 ;
#        PORT
#        LAYER M1M ;
#        RECT  3.05 4.10 3.95 5.00 ;
#        END
#    END A
#    PIN vdd!
#        DIRECTION INOUT ;
#        USE power ;
#        SHAPE ABUTMENT ;
#        PORT
#        LAYER M1M ;
#        RECT  0.45 7.15 1.15 11.00 ;
#        RECT  0.45 10.10 2.15 11.00 ;
#        RECT  3.30 7.15 4.00 11.00 ;
#        RECT  7.35 7.70 8.05 11.00 ;
#        RECT  10.05 7.70 10.75 11.00 ;
#        RECT  7.15 10.10 10.75 11.00 ;
#        RECT  0.00 11.00 11.20 13.00 ;
#        END
#    END vdd!
#    PIN gnd!
#        DIRECTION INOUT ;
#        USE ground ;
#        SHAPE ABUTMENT ;
#        PORT
#        LAYER M1M ;
#        RECT  3.50 2.00 4.20 3.65 ;
#        RECT  6.20 2.00 6.90 3.65 ;
#        RECT  10.05 2.00 10.75 3.65 ;
#        RECT  0.00 0.00 11.20 2.00 ;
#        END
#    END gnd!
#    OBS
#        LAYER M1M ;
#        RECT  0.65 2.95 1.15 6.30 ;
#        RECT  0.65 2.95 1.85 3.65 ;
#        RECT  1.80 5.80 2.50 7.85 ;
#        RECT  3.90 5.60 4.60 6.30 ;
#        RECT  0.65 5.80 4.60 6.30 ;
#        RECT  6.00 4.20 8.20 4.90 ;
#        RECT  7.70 2.95 8.20 7.25 ;
#        RECT  7.70 2.95 8.40 3.65 ;
#        RECT  7.70 6.75 9.40 7.25 ;
#        RECT  8.70 6.75 9.40 8.40 ;
#    END
#END AND4X1
MACRO AND4X2
    CLASS CORE ;
    FOREIGN AND4X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.30 4.45 5.40 4.95 ;
        RECT  4.90 2.45 5.00 7.65 ;
        RECT  4.30 2.45 5.00 4.95 ;
        RECT  4.90 4.45 5.40 7.65 ;
        RECT  4.90 7.15 6.35 7.65 ;
        RECT  5.65 7.15 6.35 9.90 ;
        RECT  5.65 8.00 6.75 9.90 ;
        RECT  5.65 9.20 9.45 9.90 ;
        RECT  8.75 9.20 9.45 10.55 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.70 1.15 11.00 ;
        RECT  0.45 10.10 2.50 11.00 ;
        RECT  3.30 7.70 4.00 11.00 ;
        RECT  7.35 7.20 8.05 8.75 ;
        RECT  7.35 8.25 10.75 8.75 ;
        RECT  10.05 7.20 10.75 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.95 2.00 3.65 4.00 ;
        RECT  5.65 2.00 6.35 4.00 ;
        RECT  10.05 2.00 10.75 4.15 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.45 1.15 4.95 ;
        RECT  1.80 6.75 2.50 8.40 ;
        RECT  0.45 4.45 3.50 4.95 ;
        RECT  3.00 4.45 3.50 7.25 ;
        RECT  1.80 6.75 3.50 7.25 ;
        RECT  3.00 5.50 4.45 6.20 ;
        RECT  5.85 4.45 6.55 5.25 ;
        RECT  7.70 3.45 8.40 4.95 ;
        RECT  5.85 4.45 9.25 4.95 ;
        RECT  8.70 4.45 9.25 7.80 ;
        RECT  8.70 7.10 9.40 7.80 ;
    END
END AND4X2
MACRO AND4X3
    CLASS CORE ;
    FOREIGN AND4X3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  5.50 9.15 10.05 9.80 ;
        RECT  7.25 2.45 8.15 4.05 ;
        RECT  7.65 2.45 8.15 7.20 ;
        RECT  7.65 6.70 9.35 7.20 ;
        RECT  8.65 6.70 9.35 9.80 ;
        RECT  5.50 9.10 9.35 9.80 ;
        RECT  9.35 9.15 10.05 10.55 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.60 1.15 11.00 ;
        RECT  0.45 10.25 2.15 11.00 ;
        RECT  3.15 6.75 3.85 11.00 ;
        RECT  3.15 6.75 7.00 7.45 ;
        RECT  10.15 7.10 11.00 8.70 ;
        RECT  10.50 7.10 11.00 11.00 ;
        RECT  12.85 7.15 13.55 11.00 ;
        RECT  10.50 10.10 13.55 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 4.05 ;
        RECT  4.45 2.00 5.15 3.95 ;
        RECT  5.95 2.00 6.65 4.00 ;
        RECT  8.65 2.00 9.35 4.00 ;
        RECT  12.50 2.00 13.20 4.05 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.00 4.50 7.20 4.95 ;
        RECT  2.00 4.45 2.50 9.30 ;
        RECT  1.80 7.60 2.50 9.30 ;
        RECT  2.80 2.45 3.50 4.95 ;
        RECT  6.50 4.45 7.00 5.20 ;
        RECT  2.00 4.45 7.00 4.95 ;
        RECT  6.50 4.50 7.20 5.20 ;
        RECT  8.60 4.45 9.30 5.25 ;
        RECT  10.15 2.45 10.85 4.95 ;
        RECT  8.60 4.45 12.05 4.95 ;
        RECT  11.50 4.45 12.05 8.85 ;
        RECT  11.50 7.15 12.20 8.85 ;
    END
END AND4X3
MACRO AND4X4
    CLASS CORE ;
    FOREIGN AND4X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.05 2.45 10.55 9.90 ;
        RECT  10.05 5.95 10.75 9.90 ;
        RECT  10.05 8.00 11.00 9.90 ;
        RECT  5.50 9.20 11.00 9.90 ;
        RECT  7.20 2.45 11.25 3.15 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.15 1.15 11.00 ;
        RECT  0.45 10.10 2.30 11.00 ;
        RECT  3.15 6.85 3.85 11.00 ;
        RECT  7.70 5.95 8.40 7.55 ;
        RECT  3.15 6.85 8.40 7.55 ;
        RECT  11.55 6.90 12.25 11.00 ;
        RECT  14.25 7.10 14.95 11.00 ;
        RECT  11.55 10.10 14.95 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 2.00 3.50 4.00 ;
        RECT  4.35 2.00 5.05 3.80 ;
        RECT  5.85 2.00 6.55 3.15 ;
        RECT  11.90 2.00 12.60 3.10 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 2.45 1.15 4.05 ;
        RECT  0.65 2.45 1.15 4.95 ;
        RECT  2.00 4.45 2.50 8.85 ;
        RECT  1.80 7.15 2.50 8.85 ;
        RECT  8.15 4.25 8.85 4.95 ;
        RECT  0.65 4.45 8.85 4.95 ;
        RECT  11.00 3.90 11.70 4.60 ;
        RECT  12.90 3.90 13.45 8.70 ;
        RECT  12.90 7.10 13.60 8.70 ;
        RECT  14.25 2.45 14.75 4.40 ;
        RECT  11.00 3.90 14.75 4.40 ;
        RECT  14.25 2.45 14.95 3.15 ;
    END
END AND4X4
MACRO AND5X1
    CLASS CORE ;
    FOREIGN AND5X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  6.25 2.95 6.95 3.65 ;
        RECT  6.45 2.95 6.95 5.90 ;
        RECT  6.45 5.40 8.15 5.90 ;
        RECT  7.05 5.40 7.75 10.55 ;
        RECT  7.05 5.40 8.15 6.30 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  11.45 4.10 12.35 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 4.10 2.55 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 3.95 5.00 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  4.45 4.10 5.35 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 7.15 2.55 11.00 ;
        RECT  0.45 10.10 3.90 11.00 ;
        RECT  4.70 7.15 5.40 11.00 ;
        RECT  8.75 7.70 9.45 11.00 ;
        RECT  11.45 7.70 12.15 11.00 ;
        RECT  8.55 10.10 12.15 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  4.90 2.00 5.60 3.65 ;
        RECT  7.60 2.00 8.30 3.65 ;
        RECT  11.45 2.00 12.15 3.65 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.70 2.95 1.20 7.85 ;
        RECT  0.50 7.15 1.20 7.85 ;
        RECT  0.70 2.95 2.20 3.65 ;
        RECT  3.20 5.80 3.90 7.85 ;
        RECT  5.30 5.60 6.00 6.30 ;
        RECT  0.70 5.80 6.00 6.30 ;
        RECT  7.40 4.20 9.60 4.90 ;
        RECT  9.10 2.95 9.60 7.25 ;
        RECT  9.10 2.95 9.80 3.65 ;
        RECT  9.10 6.75 10.80 7.25 ;
        RECT  10.10 6.75 10.80 8.40 ;
    END
END AND5X1
MACRO AND5X2
    CLASS CORE ;
    FOREIGN AND5X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  5.55 2.45 6.25 4.95 ;
        RECT  5.55 4.45 6.80 4.95 ;
        RECT  6.30 4.45 6.80 7.65 ;
        RECT  6.30 7.15 7.75 7.65 ;
        RECT  7.05 7.15 7.75 9.90 ;
        RECT  7.05 8.00 8.15 9.90 ;
        RECT  7.05 9.20 10.85 9.90 ;
        RECT  10.15 9.20 10.85 10.55 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.40 9.55 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 7.70 2.55 11.00 ;
        RECT  0.45 10.10 3.85 11.00 ;
        RECT  4.70 7.70 5.40 11.00 ;
        RECT  8.75 7.20 9.45 8.75 ;
        RECT  8.75 8.25 12.15 8.75 ;
        RECT  11.45 7.20 12.15 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  4.20 2.00 4.90 4.00 ;
        RECT  6.90 2.00 7.60 4.00 ;
        RECT  11.45 2.00 12.15 4.15 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.50 6.75 1.20 8.40 ;
        RECT  0.70 3.30 1.40 4.95 ;
        RECT  3.20 6.75 3.90 8.40 ;
        RECT  0.70 4.45 4.90 4.95 ;
        RECT  4.40 4.45 4.90 7.25 ;
        RECT  0.50 6.75 4.90 7.25 ;
        RECT  4.40 5.50 5.85 6.20 ;
        RECT  7.25 4.45 7.95 5.25 ;
        RECT  9.10 3.45 9.80 4.95 ;
        RECT  7.25 4.45 10.65 4.95 ;
        RECT  10.10 4.45 10.65 7.80 ;
        RECT  10.10 7.10 10.80 7.80 ;
    END
END AND5X2
MACRO AND5X3
    CLASS CORE ;
    FOREIGN AND5X3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  6.90 9.15 11.45 9.80 ;
        RECT  8.65 2.45 9.55 4.05 ;
        RECT  9.05 2.45 9.55 7.20 ;
        RECT  9.05 6.70 10.75 7.20 ;
        RECT  10.05 6.70 10.75 9.80 ;
        RECT  6.90 9.10 10.75 9.80 ;
        RECT  10.75 9.15 11.45 10.55 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 7.70 2.55 11.00 ;
        RECT  0.45 10.25 3.55 11.00 ;
        RECT  4.55 6.75 5.25 11.00 ;
        RECT  4.55 6.75 8.40 7.45 ;
        RECT  11.55 7.10 12.40 8.70 ;
        RECT  11.90 7.10 12.40 11.00 ;
        RECT  14.25 7.15 14.95 11.00 ;
        RECT  11.90 10.10 14.95 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.65 2.00 1.35 4.00 ;
        RECT  5.70 2.00 6.40 3.95 ;
        RECT  7.35 2.00 8.05 4.00 ;
        RECT  10.05 2.00 10.75 4.00 ;
        RECT  13.90 2.00 14.60 4.05 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.40 4.50 8.60 4.95 ;
        RECT  0.50 6.75 1.20 9.30 ;
        RECT  0.50 6.75 3.90 7.25 ;
        RECT  3.40 4.45 3.90 9.30 ;
        RECT  3.20 6.75 3.90 9.30 ;
        RECT  4.00 2.45 4.70 4.95 ;
        RECT  7.90 4.45 8.40 5.20 ;
        RECT  3.40 4.45 8.40 4.95 ;
        RECT  7.90 4.50 8.60 5.20 ;
        RECT  10.00 4.45 10.70 5.25 ;
        RECT  11.55 2.45 12.25 4.95 ;
        RECT  10.00 4.45 13.45 4.95 ;
        RECT  12.90 4.45 13.45 8.85 ;
        RECT  12.90 7.15 13.60 8.85 ;
    END
END AND5X3
MACRO AND5X4
    CLASS CORE ;
    FOREIGN AND5X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.45 2.45 11.95 9.90 ;
        RECT  11.45 5.95 12.15 9.90 ;
        RECT  11.45 8.00 12.40 9.90 ;
        RECT  6.90 9.20 12.40 9.90 ;
        RECT  8.60 2.45 12.65 3.15 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 7.70 2.55 11.00 ;
        RECT  0.45 10.20 3.75 11.00 ;
        RECT  4.55 6.85 5.25 11.00 ;
        RECT  9.10 5.95 9.80 7.55 ;
        RECT  4.55 6.85 9.80 7.55 ;
        RECT  12.95 6.90 13.65 11.00 ;
        RECT  15.65 7.10 16.35 11.00 ;
        RECT  12.95 10.10 16.35 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.85 2.00 1.55 4.00 ;
        RECT  5.75 2.00 6.45 3.80 ;
        RECT  7.25 2.00 7.95 3.15 ;
        RECT  13.30 2.00 14.00 3.10 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.50 6.75 1.20 9.25 ;
        RECT  0.50 6.75 3.90 7.25 ;
        RECT  3.40 4.45 3.90 9.25 ;
        RECT  3.20 6.75 3.90 9.25 ;
        RECT  4.20 2.45 4.90 4.95 ;
        RECT  9.55 4.25 10.25 4.95 ;
        RECT  3.40 4.45 10.25 4.95 ;
        RECT  12.40 3.90 13.10 4.60 ;
        RECT  14.30 3.90 14.85 8.70 ;
        RECT  14.30 7.10 15.00 8.70 ;
        RECT  15.65 2.45 16.15 4.40 ;
        RECT  12.40 3.90 16.15 4.40 ;
        RECT  15.65 2.45 16.35 3.15 ;
    END
END AND5X4
MACRO AND6X1
    CLASS CORE ;
    FOREIGN AND6X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  6.25 2.95 6.95 3.65 ;
        RECT  6.45 2.95 6.95 5.90 ;
        RECT  6.45 5.40 8.15 5.90 ;
        RECT  7.05 5.40 7.75 10.55 ;
        RECT  7.05 5.40 8.15 6.30 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 4.10 2.55 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 3.95 5.00 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  4.45 4.10 5.35 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 7.15 2.55 11.00 ;
        RECT  0.45 10.10 3.90 11.00 ;
        RECT  4.70 7.15 5.40 11.00 ;
        RECT  8.75 7.70 9.45 11.00 ;
        RECT  11.45 7.70 12.15 11.00 ;
        RECT  8.75 10.10 13.55 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  4.90 2.00 5.60 3.65 ;
        RECT  7.60 2.00 8.30 3.65 ;
        RECT  12.80 2.00 13.50 3.90 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.70 2.70 1.20 7.85 ;
        RECT  0.50 7.15 1.20 7.85 ;
        RECT  0.70 2.70 2.20 3.40 ;
        RECT  3.20 5.80 3.90 7.85 ;
        RECT  5.30 5.60 6.00 6.30 ;
        RECT  0.70 5.80 6.00 6.30 ;
        RECT  7.40 4.20 9.60 4.90 ;
        RECT  9.10 3.20 9.60 7.25 ;
        RECT  9.10 3.20 10.15 3.90 ;
        RECT  10.10 6.75 10.80 8.40 ;
        RECT  9.10 6.75 13.50 7.25 ;
        RECT  12.80 6.75 13.50 8.40 ;
    END
END AND6X1
MACRO AND6X2
    CLASS CORE ;
    FOREIGN AND6X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  5.35 2.45 6.05 4.95 ;
        RECT  5.35 4.45 6.60 4.95 ;
        RECT  6.10 4.45 6.60 7.65 ;
        RECT  6.10 7.15 7.70 7.65 ;
        RECT  7.25 7.15 7.70 10.20 ;
        RECT  7.00 7.15 7.70 9.90 ;
        RECT  7.25 9.20 8.15 10.20 ;
        RECT  7.00 9.20 10.80 9.90 ;
        RECT  10.10 9.20 10.80 10.50 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.40 9.55 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.70 2.50 11.00 ;
        RECT  0.45 10.10 3.85 11.00 ;
        RECT  4.65 7.70 5.35 11.00 ;
        RECT  8.50 7.70 9.20 8.75 ;
        RECT  8.50 8.25 12.20 8.75 ;
        RECT  11.50 7.70 12.20 11.00 ;
        RECT  11.50 10.10 13.45 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  4.00 2.00 4.70 4.00 ;
        RECT  6.70 2.00 7.40 4.00 ;
        RECT  12.50 2.00 13.20 4.15 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 6.75 1.15 8.40 ;
        RECT  0.50 3.25 1.20 4.95 ;
        RECT  3.15 6.75 3.85 8.40 ;
        RECT  0.50 4.45 4.90 4.95 ;
        RECT  4.40 4.45 4.90 7.25 ;
        RECT  0.45 6.75 4.90 7.25 ;
        RECT  4.40 5.50 5.65 6.20 ;
        RECT  7.05 4.45 7.75 5.25 ;
        RECT  9.15 3.45 9.85 4.95 ;
        RECT  7.05 4.45 10.50 4.95 ;
        RECT  10.00 4.45 10.50 7.80 ;
        RECT  10.00 6.75 10.70 7.80 ;
        RECT  10.00 6.75 13.55 7.25 ;
        RECT  12.85 6.75 13.55 8.40 ;
    END
END AND6X2
MACRO AND6X3
    CLASS CORE ;
    FOREIGN AND6X3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  6.90 9.15 11.45 9.80 ;
        RECT  8.15 2.45 8.85 4.05 ;
        RECT  8.35 2.45 8.85 6.30 ;
        RECT  8.35 5.80 10.75 6.30 ;
        RECT  10.05 5.80 10.75 9.80 ;
        RECT  10.75 8.00 10.95 10.55 ;
        RECT  6.90 9.10 10.95 9.80 ;
        RECT  10.75 9.15 11.45 10.55 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 7.70 2.55 11.00 ;
        RECT  0.45 10.25 3.55 11.00 ;
        RECT  4.55 6.75 5.25 11.00 ;
        RECT  4.55 6.75 8.40 7.45 ;
        RECT  11.55 7.10 12.40 8.70 ;
        RECT  11.90 7.10 12.40 11.00 ;
        RECT  14.25 7.70 14.95 11.00 ;
        RECT  11.90 10.10 16.30 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 4.00 ;
        RECT  5.30 2.00 6.00 3.95 ;
        RECT  6.80 2.00 7.50 4.00 ;
        RECT  9.50 2.00 10.20 4.00 ;
        RECT  15.65 2.00 16.35 4.00 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.50 6.75 1.20 9.30 ;
        RECT  0.50 6.75 3.90 7.25 ;
        RECT  3.40 4.45 3.90 9.30 ;
        RECT  3.80 2.45 3.90 9.30 ;
        RECT  3.20 6.75 3.90 9.30 ;
        RECT  3.80 2.45 4.50 4.95 ;
        RECT  3.40 4.45 7.80 4.95 ;
        RECT  7.10 4.45 7.80 5.15 ;
        RECT  9.30 4.45 10.00 5.25 ;
        RECT  9.30 4.45 13.45 4.95 ;
        RECT  12.90 2.45 13.00 8.85 ;
        RECT  12.30 2.45 13.00 4.95 ;
        RECT  12.90 4.45 13.45 8.85 ;
        RECT  12.90 6.75 13.60 8.85 ;
        RECT  12.90 6.75 16.30 7.25 ;
        RECT  15.60 6.75 16.30 9.05 ;
    END
END AND6X3
MACRO AND6X4
    CLASS CORE ;
    FOREIGN AND6X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  9.20 2.45 9.90 4.05 ;
        RECT  9.20 2.45 11.45 3.15 ;
        RECT  10.75 2.45 11.25 6.30 ;
        RECT  10.75 2.45 11.45 4.05 ;
        RECT  10.75 5.80 13.40 6.30 ;
        RECT  6.90 9.20 13.40 9.90 ;
        RECT  12.70 5.80 13.40 10.55 ;
        RECT  12.70 8.00 13.75 8.90 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.40 19.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 7.75 2.55 11.00 ;
        RECT  0.50 10.35 3.70 11.00 ;
        RECT  4.55 6.85 5.25 11.00 ;
        RECT  4.55 6.85 10.85 7.55 ;
        RECT  14.20 7.60 14.90 11.00 ;
        RECT  17.05 7.70 17.75 11.00 ;
        RECT  14.20 10.20 19.15 11.00 ;
        RECT  0.00 11.00 19.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 4.40 ;
        RECT  5.40 2.00 7.00 3.80 ;
        RECT  7.85 2.00 8.55 4.00 ;
        RECT  12.10 2.00 12.80 4.00 ;
        RECT  13.60 2.00 14.30 3.80 ;
        RECT  18.45 2.00 19.15 4.40 ;
        RECT  0.00 0.00 19.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.50 6.80 1.20 9.35 ;
        RECT  0.50 6.80 3.90 7.30 ;
        RECT  3.40 4.45 3.90 9.35 ;
        RECT  3.80 2.45 3.90 9.35 ;
        RECT  3.20 6.80 3.90 9.35 ;
        RECT  3.80 2.45 4.50 4.95 ;
        RECT  3.40 4.45 8.95 4.95 ;
        RECT  8.25 4.45 8.95 5.15 ;
        RECT  11.70 4.45 12.40 5.15 ;
        RECT  11.70 4.45 16.25 4.95 ;
        RECT  15.75 2.45 15.80 9.25 ;
        RECT  15.10 2.45 15.80 4.95 ;
        RECT  15.75 4.45 16.25 9.25 ;
        RECT  15.55 6.75 16.25 9.25 ;
        RECT  15.55 6.75 19.10 7.25 ;
        RECT  18.40 6.75 19.10 9.25 ;
    END
END AND6X4
MACRO AND7X1
    CLASS CORE ;
    FOREIGN AND7X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  6.25 3.00 6.95 4.60 ;
        RECT  7.05 4.10 7.55 6.95 ;
        RECT  7.05 6.45 9.15 6.95 ;
        RECT  8.45 6.45 9.15 10.55 ;
        RECT  8.45 8.00 9.55 8.90 ;
        RECT  8.95 3.00 9.65 4.60 ;
        RECT  6.25 4.10 9.65 4.60 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  14.25 9.30 15.15 10.20 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  4.45 4.10 5.35 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 3.95 5.00 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 4.10 2.55 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.20 7.15 2.90 11.00 ;
        RECT  0.45 10.10 3.90 11.00 ;
        RECT  5.10 6.65 5.80 11.00 ;
        RECT  10.25 7.70 10.95 11.00 ;
        RECT  12.95 7.70 13.65 11.00 ;
        RECT  9.95 10.10 13.65 11.00 ;
        RECT  15.65 7.70 16.35 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  4.90 2.00 5.60 3.65 ;
        RECT  7.60 2.00 8.30 3.65 ;
        RECT  12.95 2.00 13.65 4.30 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.85 2.70 1.20 7.85 ;
        RECT  0.70 2.70 1.20 6.00 ;
        RECT  0.85 5.50 1.55 7.85 ;
        RECT  0.70 2.70 2.20 3.40 ;
        RECT  3.55 5.50 4.25 7.85 ;
        RECT  5.70 5.30 6.40 6.00 ;
        RECT  0.70 5.50 6.40 6.00 ;
        RECT  8.00 5.30 8.70 6.00 ;
        RECT  8.00 5.30 10.95 5.80 ;
        RECT  10.45 2.75 10.95 7.25 ;
        RECT  10.45 2.75 11.15 3.45 ;
        RECT  10.45 6.75 12.30 7.25 ;
        RECT  11.60 6.75 12.30 8.40 ;
        RECT  14.50 3.75 15.00 8.40 ;
        RECT  14.30 7.70 15.00 8.40 ;
        RECT  15.45 2.45 16.15 4.25 ;
        RECT  14.50 3.75 16.15 4.25 ;
        RECT  15.45 2.45 16.50 3.15 ;
    END
END AND7X1
MACRO AND7X2
    CLASS CORE ;
    FOREIGN AND7X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  7.50 3.00 8.20 4.60 ;
        RECT  10.20 3.00 10.90 4.60 ;
        RECT  12.90 3.00 13.60 4.60 ;
        RECT  7.50 4.10 14.90 4.60 ;
        RECT  14.25 8.00 15.15 8.90 ;
        RECT  14.40 4.10 14.90 9.60 ;
        RECT  14.40 6.60 15.15 9.60 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.40 19.35 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  17.05 4.10 17.95 5.00 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  19.85 4.10 20.75 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  22.65 5.40 23.55 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.70 2.50 11.00 ;
        RECT  0.50 10.10 3.65 11.00 ;
        RECT  4.65 7.70 5.35 11.00 ;
        RECT  7.35 7.40 8.05 11.00 ;
        RECT  17.25 7.70 17.95 11.00 ;
        RECT  19.95 7.70 20.65 11.00 ;
        RECT  22.65 7.70 23.35 11.00 ;
        RECT  17.25 10.10 23.35 11.00 ;
        RECT  0.00 11.00 23.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.65 ;
        RECT  6.15 2.00 6.85 3.65 ;
        RECT  8.85 2.00 9.55 3.65 ;
        RECT  11.55 2.00 12.25 3.65 ;
        RECT  14.25 2.00 14.95 3.65 ;
        RECT  19.40 2.00 20.10 3.65 ;
        RECT  0.00 0.00 23.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 6.75 1.15 8.40 ;
        RECT  3.15 6.75 3.85 8.40 ;
        RECT  3.80 2.70 4.90 3.40 ;
        RECT  4.40 2.70 4.90 7.25 ;
        RECT  0.45 6.75 4.90 7.25 ;
        RECT  4.40 5.30 6.25 6.00 ;
        RECT  6.00 6.45 6.70 10.55 ;
        RECT  6.00 6.45 9.55 6.95 ;
        RECT  8.85 6.45 9.55 10.55 ;
        RECT  10.20 6.45 10.90 9.60 ;
        RECT  11.55 7.40 12.25 10.55 ;
        RECT  8.85 10.05 12.25 10.55 ;
        RECT  10.20 6.45 13.75 6.95 ;
        RECT  13.05 6.45 13.75 10.55 ;
        RECT  15.75 6.45 16.45 10.55 ;
        RECT  13.05 10.05 16.45 10.55 ;
        RECT  16.10 2.95 16.60 6.00 ;
        RECT  15.35 5.30 16.60 6.00 ;
        RECT  15.35 5.50 17.75 6.00 ;
        RECT  16.10 2.95 17.75 3.65 ;
        RECT  17.25 5.50 17.75 7.25 ;
        RECT  17.25 6.75 19.30 7.25 ;
        RECT  18.60 6.75 19.30 8.40 ;
        RECT  21.50 3.00 22.00 8.40 ;
        RECT  21.30 7.70 22.00 8.40 ;
        RECT  22.80 2.45 23.50 3.70 ;
        RECT  21.50 3.00 23.50 3.70 ;
    END
END AND7X2
MACRO AND7X3
    CLASS CORE ;
    FOREIGN AND7X3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 25.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.70 4.10 15.15 4.35 ;
        RECT  8.70 2.75 9.40 4.35 ;
        RECT  11.40 2.75 12.10 4.35 ;
        RECT  14.10 2.75 14.60 9.60 ;
        RECT  14.10 2.75 14.80 5.00 ;
        RECT  8.70 3.85 14.80 4.35 ;
        RECT  14.10 6.45 14.80 9.60 ;
        RECT  14.10 4.10 15.15 5.00 ;
        RECT  14.10 6.45 17.50 6.95 ;
        RECT  16.80 6.45 17.50 10.55 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  18.45 4.10 19.35 5.00 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  21.25 4.10 22.15 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  24.05 5.40 24.95 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.70 2.50 11.00 ;
        RECT  0.50 10.35 3.65 11.00 ;
        RECT  4.65 7.70 5.35 11.00 ;
        RECT  7.35 7.40 8.05 11.00 ;
        RECT  18.65 7.70 19.35 11.00 ;
        RECT  21.35 7.70 22.05 11.00 ;
        RECT  24.05 7.70 24.75 11.00 ;
        RECT  18.65 10.35 24.75 11.00 ;
        RECT  0.00 11.00 25.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.95 2.00 4.65 3.65 ;
        RECT  5.50 2.00 6.20 3.80 ;
        RECT  7.35 2.00 8.05 3.40 ;
        RECT  10.05 2.00 10.75 3.40 ;
        RECT  12.75 2.00 13.45 3.40 ;
        RECT  15.45 2.00 16.15 3.40 ;
        RECT  20.80 2.00 21.50 3.65 ;
        RECT  0.00 0.00 25.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 2.45 1.15 4.60 ;
        RECT  0.45 6.75 1.15 9.40 ;
        RECT  3.15 6.75 3.85 9.40 ;
        RECT  0.45 4.10 4.90 4.60 ;
        RECT  4.40 4.10 4.90 7.25 ;
        RECT  0.45 6.75 4.90 7.25 ;
        RECT  4.40 5.30 6.25 6.00 ;
        RECT  6.00 6.45 6.70 10.55 ;
        RECT  6.00 6.45 9.40 6.95 ;
        RECT  8.70 6.45 9.40 10.55 ;
        RECT  10.05 6.45 10.75 9.60 ;
        RECT  11.40 7.40 12.10 10.55 ;
        RECT  8.70 10.05 12.10 10.55 ;
        RECT  10.05 6.45 13.45 6.95 ;
        RECT  12.75 6.45 13.45 10.55 ;
        RECT  15.45 7.40 16.15 10.55 ;
        RECT  12.75 10.05 16.15 10.55 ;
        RECT  15.90 5.30 16.60 6.00 ;
        RECT  15.90 5.50 18.50 6.00 ;
        RECT  17.50 2.50 18.00 6.00 ;
        RECT  18.00 5.50 18.50 7.25 ;
        RECT  17.50 2.50 19.15 3.20 ;
        RECT  18.00 6.75 20.70 7.25 ;
        RECT  20.00 6.75 20.70 9.40 ;
        RECT  22.90 2.45 23.40 9.40 ;
        RECT  22.70 7.70 23.40 9.40 ;
        RECT  22.90 2.45 24.90 3.25 ;
    END
END AND7X3
MACRO AND7X4
    CLASS CORE ;
    FOREIGN AND7X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 32.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.55 2.50 12.25 4.70 ;
        RECT  14.25 2.50 14.95 4.70 ;
        RECT  16.95 2.50 17.65 4.70 ;
        RECT  11.55 4.20 20.30 4.70 ;
        RECT  19.80 4.20 20.30 9.60 ;
        RECT  19.80 5.40 20.50 9.60 ;
        RECT  19.80 5.40 20.75 6.95 ;
        RECT  19.80 6.45 23.20 6.95 ;
        RECT  22.50 6.45 23.20 9.60 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  26.85 5.40 27.75 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  25.45 5.40 26.35 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  31.05 5.40 31.95 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  28.25 4.10 29.15 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.70 2.50 11.00 ;
        RECT  0.50 10.35 3.65 11.00 ;
        RECT  4.65 7.70 5.35 11.00 ;
        RECT  7.35 7.40 8.05 11.00 ;
        RECT  10.05 7.40 10.75 11.00 ;
        RECT  25.35 7.70 26.05 11.00 ;
        RECT  28.05 7.70 28.75 11.00 ;
        RECT  30.75 7.70 31.45 11.00 ;
        RECT  25.35 10.35 31.75 11.00 ;
        RECT  0.00 11.00 32.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.95 2.00 4.65 3.65 ;
        RECT  5.95 2.00 9.35 3.80 ;
        RECT  10.20 2.00 10.90 3.65 ;
        RECT  12.90 2.00 13.60 3.65 ;
        RECT  15.60 2.00 16.30 3.65 ;
        RECT  18.30 2.00 19.00 3.65 ;
        RECT  19.80 2.00 23.20 3.75 ;
        RECT  26.50 2.00 27.20 3.65 ;
        RECT  31.05 2.00 31.75 3.75 ;
        RECT  0.00 0.00 32.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 2.45 1.15 4.60 ;
        RECT  0.45 6.75 1.15 9.40 ;
        RECT  3.15 6.75 3.85 9.40 ;
        RECT  0.45 4.10 4.90 4.60 ;
        RECT  4.40 4.10 4.90 7.25 ;
        RECT  0.45 6.75 4.90 7.25 ;
        RECT  4.40 5.30 6.25 6.00 ;
        RECT  6.00 6.45 6.70 10.55 ;
        RECT  8.70 6.45 9.40 10.55 ;
        RECT  6.00 6.45 12.25 6.95 ;
        RECT  11.55 6.45 12.25 10.55 ;
        RECT  12.90 6.45 13.60 9.60 ;
        RECT  14.25 7.40 14.95 10.55 ;
        RECT  15.60 6.45 16.30 9.60 ;
        RECT  16.95 7.40 17.65 10.55 ;
        RECT  11.55 10.05 17.65 10.55 ;
        RECT  12.90 6.45 19.15 6.95 ;
        RECT  18.45 6.45 19.15 10.55 ;
        RECT  21.15 7.40 21.85 10.55 ;
        RECT  22.95 5.30 24.65 6.00 ;
        RECT  23.85 7.70 24.55 10.55 ;
        RECT  18.45 10.05 24.55 10.55 ;
        RECT  24.15 2.50 24.65 7.25 ;
        RECT  24.15 2.50 24.85 3.20 ;
        RECT  24.15 6.75 27.40 7.25 ;
        RECT  26.70 6.75 27.40 9.40 ;
        RECT  27.65 2.55 30.15 3.30 ;
        RECT  29.65 2.55 30.15 9.40 ;
        RECT  29.40 7.70 30.15 9.40 ;
    END
END AND7X4
MACRO AND8X1
    CLASS CORE ;
    FOREIGN AND8X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  6.25 3.00 6.95 4.60 ;
        RECT  7.05 4.10 7.55 6.95 ;
        RECT  7.05 6.45 9.15 6.95 ;
        RECT  8.45 6.45 9.15 10.55 ;
        RECT  8.45 8.00 9.55 8.90 ;
        RECT  8.95 3.00 9.65 4.60 ;
        RECT  6.25 4.10 9.65 4.60 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  15.65 9.30 16.55 10.20 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  4.45 4.10 5.35 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 3.95 5.00 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 4.10 2.55 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.20 7.15 2.90 11.00 ;
        RECT  0.45 10.10 3.90 11.00 ;
        RECT  5.10 6.65 5.80 11.00 ;
        RECT  11.65 7.70 12.35 11.00 ;
        RECT  14.35 7.70 15.05 11.00 ;
        RECT  9.95 10.10 15.05 11.00 ;
        RECT  17.05 7.70 17.75 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  4.90 2.00 5.60 3.65 ;
        RECT  7.60 2.00 8.30 3.65 ;
        RECT  14.35 2.00 15.05 4.00 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.85 2.70 1.20 7.85 ;
        RECT  0.70 2.70 1.20 6.00 ;
        RECT  0.85 5.50 1.55 7.85 ;
        RECT  0.70 2.70 2.20 3.40 ;
        RECT  3.55 5.50 4.25 7.85 ;
        RECT  5.70 5.30 6.40 6.00 ;
        RECT  0.70 5.50 6.40 6.00 ;
        RECT  8.00 5.30 8.70 6.00 ;
        RECT  8.00 5.30 11.00 5.80 ;
        RECT  10.50 3.05 11.00 8.40 ;
        RECT  10.30 6.75 11.00 8.40 ;
        RECT  10.50 3.05 11.70 3.75 ;
        RECT  10.30 6.75 13.70 7.25 ;
        RECT  13.00 6.75 13.70 8.40 ;
        RECT  15.90 3.75 16.40 8.40 ;
        RECT  15.70 7.70 16.40 8.40 ;
        RECT  16.85 2.45 17.55 4.25 ;
        RECT  15.90 3.75 17.55 4.25 ;
        RECT  16.85 2.45 17.90 3.15 ;
    END
END AND8X1
MACRO AND8X2
    CLASS CORE ;
    FOREIGN AND8X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 25.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  7.50 3.00 8.20 4.60 ;
        RECT  10.20 3.00 10.90 4.60 ;
        RECT  12.90 3.00 13.60 4.60 ;
        RECT  7.50 4.10 14.90 4.60 ;
        RECT  14.25 8.00 15.15 8.90 ;
        RECT  14.40 4.10 14.90 9.60 ;
        RECT  14.40 6.60 15.15 9.60 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.40 19.35 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  21.25 4.10 22.15 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  24.05 5.40 24.95 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.70 2.50 11.00 ;
        RECT  0.50 10.10 3.65 11.00 ;
        RECT  4.65 7.70 5.35 11.00 ;
        RECT  7.35 7.40 8.05 11.00 ;
        RECT  18.65 7.70 19.35 11.00 ;
        RECT  21.35 7.70 22.05 11.00 ;
        RECT  24.05 7.70 24.75 11.00 ;
        RECT  17.55 10.10 24.75 11.00 ;
        RECT  0.00 11.00 25.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.45 ;
        RECT  6.15 2.00 6.85 3.65 ;
        RECT  8.85 2.00 9.55 3.65 ;
        RECT  11.55 2.00 12.25 3.65 ;
        RECT  14.25 2.00 14.95 3.65 ;
        RECT  20.80 2.00 21.50 3.65 ;
        RECT  0.00 0.00 25.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 6.75 1.15 8.40 ;
        RECT  3.15 6.75 3.85 8.40 ;
        RECT  3.80 2.75 4.90 3.45 ;
        RECT  4.40 2.75 4.90 7.25 ;
        RECT  0.45 6.75 4.90 7.25 ;
        RECT  4.40 5.30 6.25 6.00 ;
        RECT  6.00 6.45 6.70 10.55 ;
        RECT  6.00 6.45 9.55 6.95 ;
        RECT  8.85 6.45 9.55 10.55 ;
        RECT  10.20 6.45 10.90 9.60 ;
        RECT  11.55 7.40 12.25 10.55 ;
        RECT  8.85 10.05 12.25 10.55 ;
        RECT  10.20 6.45 13.75 6.95 ;
        RECT  13.05 6.45 13.75 10.55 ;
        RECT  15.35 5.30 16.60 6.00 ;
        RECT  15.75 7.70 16.45 10.55 ;
        RECT  13.05 10.05 16.45 10.55 ;
        RECT  16.10 2.75 16.60 7.25 ;
        RECT  17.30 6.75 18.00 8.40 ;
        RECT  16.10 2.75 18.15 3.45 ;
        RECT  16.10 6.75 20.70 7.25 ;
        RECT  20.00 6.75 20.70 8.40 ;
        RECT  22.90 3.00 23.40 8.40 ;
        RECT  22.70 7.70 23.40 8.40 ;
        RECT  24.20 2.45 24.90 3.70 ;
        RECT  22.90 3.00 24.90 3.70 ;
    END
END AND8X2
MACRO AND8X3
    CLASS CORE ;
    FOREIGN AND8X3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 26.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  7.35 2.75 8.05 4.40 ;
        RECT  10.05 2.75 10.75 4.40 ;
        RECT  12.75 2.75 13.45 4.40 ;
        RECT  7.35 3.90 15.15 4.40 ;
        RECT  14.10 3.90 14.60 9.60 ;
        RECT  14.10 6.75 14.80 9.60 ;
        RECT  14.10 3.90 15.15 5.05 ;
        RECT  14.10 6.75 17.50 7.25 ;
        RECT  16.80 6.75 17.50 10.55 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  25.45 5.40 26.35 6.30 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  24.05 5.40 24.95 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  21.25 5.40 22.15 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  19.85 4.10 20.75 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  18.45 4.10 19.35 5.35 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.70 2.50 11.00 ;
        RECT  0.50 10.35 3.65 11.00 ;
        RECT  4.65 7.70 5.35 11.00 ;
        RECT  7.35 7.40 8.05 11.00 ;
        RECT  18.35 7.70 19.05 11.00 ;
        RECT  21.05 7.70 21.75 11.00 ;
        RECT  23.75 7.70 24.45 11.00 ;
        RECT  18.35 10.35 26.15 11.00 ;
        RECT  0.00 11.00 26.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.95 2.00 4.65 3.65 ;
        RECT  6.00 2.00 6.70 3.45 ;
        RECT  8.70 2.00 9.40 3.45 ;
        RECT  11.40 2.00 12.10 3.45 ;
        RECT  14.10 2.00 14.80 3.45 ;
        RECT  19.90 2.00 20.60 3.40 ;
        RECT  25.45 2.00 26.15 3.95 ;
        RECT  0.00 0.00 26.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  22.10 3.35 23.10 4.05 ;
        RECT  0.45 2.45 1.15 4.60 ;
        RECT  0.45 6.75 1.15 9.40 ;
        RECT  3.15 6.75 3.85 9.40 ;
        RECT  0.45 4.10 4.90 4.60 ;
        RECT  4.40 4.10 4.90 7.25 ;
        RECT  0.45 6.75 4.90 7.25 ;
        RECT  4.40 5.30 6.25 6.00 ;
        RECT  6.00 6.45 6.70 10.55 ;
        RECT  6.00 6.45 9.40 6.95 ;
        RECT  8.70 6.45 9.40 10.55 ;
        RECT  10.05 6.45 10.75 9.60 ;
        RECT  11.40 7.40 12.10 10.55 ;
        RECT  8.70 10.05 12.10 10.55 ;
        RECT  10.05 6.45 13.45 6.95 ;
        RECT  12.75 6.45 13.45 10.55 ;
        RECT  15.25 2.50 15.95 3.20 ;
        RECT  15.45 7.70 16.15 10.55 ;
        RECT  12.75 10.05 16.15 10.55 ;
        RECT  15.25 2.50 18.25 3.00 ;
        RECT  17.50 2.50 18.00 6.30 ;
        RECT  17.50 2.50 18.25 3.20 ;
        RECT  17.50 5.80 20.40 6.30 ;
        RECT  19.70 5.80 20.40 9.40 ;
        RECT  21.05 2.45 22.80 3.15 ;
        RECT  22.60 2.45 22.80 9.40 ;
        RECT  22.10 2.45 22.80 4.05 ;
        RECT  22.60 3.35 23.10 9.40 ;
        RECT  22.40 6.75 23.15 9.40 ;
        RECT  22.40 6.75 25.80 7.25 ;
        RECT  25.10 6.75 25.80 9.40 ;
    END
END AND8X3
MACRO AND8X4
    CLASS CORE ;
    FOREIGN AND8X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 33.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  12.90 2.50 13.60 4.70 ;
        RECT  15.60 2.50 16.30 4.70 ;
        RECT  18.30 2.50 19.00 4.70 ;
        RECT  12.90 4.20 20.30 4.70 ;
        RECT  19.80 4.20 20.30 9.60 ;
        RECT  19.80 5.40 20.50 9.60 ;
        RECT  19.80 5.40 20.75 6.95 ;
        RECT  19.80 6.45 23.20 6.95 ;
        RECT  22.50 6.45 23.20 9.60 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  32.45 5.40 33.35 6.30 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  31.05 5.40 31.95 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  28.25 5.40 29.15 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  26.85 5.40 27.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  25.45 5.40 26.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.70 2.50 11.00 ;
        RECT  0.50 10.35 3.65 11.00 ;
        RECT  4.65 7.70 5.35 11.00 ;
        RECT  7.35 7.40 8.05 11.00 ;
        RECT  10.05 7.40 10.75 11.00 ;
        RECT  25.35 7.70 26.05 11.00 ;
        RECT  28.05 7.70 28.75 11.00 ;
        RECT  30.75 7.70 31.45 11.00 ;
        RECT  25.35 10.35 33.15 11.00 ;
        RECT  0.00 11.00 33.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.95 2.00 4.65 3.65 ;
        RECT  5.50 2.00 10.70 3.80 ;
        RECT  11.55 2.00 12.25 3.65 ;
        RECT  14.25 2.00 14.95 3.65 ;
        RECT  16.95 2.00 17.65 3.65 ;
        RECT  19.65 2.00 20.35 3.65 ;
        RECT  22.35 2.00 23.05 3.80 ;
        RECT  26.90 2.00 27.60 3.65 ;
        RECT  32.45 2.00 33.15 3.95 ;
        RECT  0.00 0.00 33.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  29.10 3.35 30.10 4.05 ;
        RECT  0.45 2.45 1.15 4.60 ;
        RECT  0.45 6.75 1.15 9.40 ;
        RECT  3.15 6.75 3.85 9.40 ;
        RECT  0.45 4.10 4.90 4.60 ;
        RECT  4.40 4.10 4.90 7.25 ;
        RECT  0.45 6.75 4.90 7.25 ;
        RECT  4.40 5.30 6.25 6.00 ;
        RECT  6.00 6.45 6.70 10.55 ;
        RECT  8.70 6.45 9.40 10.55 ;
        RECT  6.00 6.45 12.25 6.95 ;
        RECT  11.55 6.45 12.25 10.55 ;
        RECT  12.90 6.45 13.60 9.60 ;
        RECT  14.25 7.40 14.95 10.55 ;
        RECT  15.60 6.45 16.30 9.60 ;
        RECT  16.95 7.40 17.65 10.55 ;
        RECT  11.55 10.05 17.65 10.55 ;
        RECT  12.90 6.45 19.15 6.95 ;
        RECT  18.45 6.45 19.15 10.55 ;
        RECT  20.80 2.45 21.50 3.15 ;
        RECT  21.00 2.45 21.50 4.85 ;
        RECT  21.15 7.40 21.85 10.55 ;
        RECT  21.00 4.35 25.00 4.85 ;
        RECT  23.85 7.70 24.55 10.55 ;
        RECT  18.45 10.05 24.55 10.55 ;
        RECT  24.50 2.50 25.00 7.25 ;
        RECT  24.50 2.50 25.25 3.20 ;
        RECT  24.50 6.75 27.40 7.25 ;
        RECT  26.70 6.75 27.40 9.40 ;
        RECT  28.05 2.45 29.80 3.15 ;
        RECT  29.60 2.45 29.80 9.40 ;
        RECT  29.10 2.45 29.80 4.05 ;
        RECT  29.60 3.35 30.10 9.40 ;
        RECT  29.40 6.75 30.15 9.40 ;
        RECT  29.40 6.75 32.80 7.25 ;
        RECT  32.10 6.75 32.80 9.40 ;
    END
END AND8X4
MACRO ANTENNACELL
    CLASS CORE FEEDTHRU ;
    FOREIGN ANTENNACELL 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 1.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.25 8.00 1.15 8.90 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.00 11.00 1.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.00 0.00 1.40 2.00 ;
        END
    END gnd!
END ANTENNACELL
MACRO AO211X1
    CLASS CORE ;
    FOREIGN AO211X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.65 3.00 9.40 3.70 ;
        RECT  8.90 3.00 9.40 8.90 ;
        RECT  8.65 7.15 9.40 8.90 ;
        RECT  8.65 8.00 9.55 8.90 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  5.85 4.10 6.75 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 3.95 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.35 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.15 7.70 2.85 11.00 ;
        RECT  7.35 7.15 8.05 11.00 ;
        RECT  7.35 10.10 10.75 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.65 ;
        RECT  4.30 2.00 5.00 2.70 ;
        RECT  7.30 2.00 8.00 3.70 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.80 6.75 1.50 10.55 ;
        RECT  0.80 6.75 4.20 7.25 ;
        RECT  2.80 2.45 3.50 3.65 ;
        RECT  3.50 6.75 4.20 10.55 ;
        RECT  4.60 3.15 5.10 6.00 ;
        RECT  5.80 2.45 6.50 3.65 ;
        RECT  2.80 3.15 6.50 3.65 ;
        RECT  5.85 5.50 6.55 10.55 ;
        RECT  7.75 5.30 8.45 6.00 ;
        RECT  4.60 5.50 8.45 6.00 ;
    END
END AO211X1
MACRO AO211X2
    CLASS CORE ;
    FOREIGN AO211X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.85 2.45 9.40 10.55 ;
        RECT  8.65 7.15 9.40 10.55 ;
        RECT  8.85 2.45 9.55 4.05 ;
        RECT  8.65 8.00 9.55 10.55 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  5.85 4.10 6.75 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 3.95 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.35 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.15 7.70 2.85 11.00 ;
        RECT  7.35 7.15 8.05 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.65 ;
        RECT  4.30 2.00 5.00 2.70 ;
        RECT  7.30 2.00 8.00 3.70 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.80 6.75 1.50 10.55 ;
        RECT  0.80 6.75 4.20 7.25 ;
        RECT  2.80 2.45 3.50 3.65 ;
        RECT  3.50 6.75 4.20 10.55 ;
        RECT  4.60 3.15 5.10 6.00 ;
        RECT  5.80 2.45 6.50 3.65 ;
        RECT  2.80 3.15 6.50 3.65 ;
        RECT  5.85 5.50 6.55 10.55 ;
        RECT  7.70 5.30 8.40 6.00 ;
        RECT  4.60 5.50 8.40 6.00 ;
    END
END AO211X2
MACRO AO211X4
    CLASS CORE ;
    FOREIGN AO211X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.70 2.50 9.40 4.10 ;
        RECT  8.85 2.50 9.40 10.55 ;
        RECT  8.65 7.15 9.40 10.55 ;
        RECT  8.65 8.00 9.55 10.55 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  5.85 4.10 6.75 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 3.95 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.35 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.15 7.70 2.85 11.00 ;
        RECT  7.35 7.15 8.05 11.00 ;
        RECT  10.05 7.15 10.75 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.65 ;
        RECT  4.30 2.00 5.00 2.70 ;
        RECT  10.05 2.00 10.75 4.40 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.80 6.75 1.50 10.55 ;
        RECT  0.80 6.75 4.20 7.25 ;
        RECT  2.80 2.45 3.50 3.65 ;
        RECT  3.50 6.75 4.20 10.55 ;
        RECT  4.75 3.15 5.25 6.00 ;
        RECT  5.80 2.45 6.50 3.65 ;
        RECT  2.80 3.15 6.50 3.65 ;
        RECT  5.85 5.50 6.55 10.55 ;
        RECT  7.70 5.30 8.40 6.00 ;
        RECT  4.75 5.50 8.40 6.00 ;
    END
END AO211X4
MACRO AO21X1
    CLASS CORE ;
    FOREIGN AO21X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.65 4.90 0.75 9.05 ;
        RECT  0.25 5.40 0.75 9.05 ;
        RECT  0.25 8.55 1.80 9.05 ;
        RECT  0.65 4.90 1.15 6.30 ;
        RECT  0.25 5.40 1.15 6.30 ;
        RECT  1.10 8.55 1.80 9.25 ;
        RECT  0.65 4.90 2.55 5.40 ;
        RECT  2.05 2.75 2.55 5.40 ;
        RECT  2.05 2.75 2.75 3.45 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 3.95 5.35 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  5.45 5.40 6.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.20 7.20 1.90 7.90 ;
        RECT  1.20 7.40 2.75 7.90 ;
        RECT  2.25 7.40 2.75 11.00 ;
        RECT  1.20 9.90 2.75 11.00 ;
        RECT  5.90 7.80 6.60 11.00 ;
        RECT  0.00 11.00 8.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 4.45 ;
        RECT  3.40 2.00 4.10 3.45 ;
        RECT  7.25 2.00 7.95 4.50 ;
        RECT  0.00 0.00 8.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.40 5.85 3.70 6.60 ;
        RECT  3.20 5.85 3.70 10.55 ;
        RECT  3.20 7.20 3.90 10.55 ;
        RECT  4.45 4.00 4.95 6.35 ;
        RECT  4.90 2.70 4.95 6.35 ;
        RECT  2.40 5.85 4.95 6.35 ;
        RECT  4.55 6.80 5.25 10.55 ;
        RECT  4.90 2.70 5.60 4.50 ;
        RECT  4.45 4.00 5.60 4.50 ;
        RECT  4.55 6.80 7.95 7.30 ;
        RECT  7.25 6.80 7.95 10.55 ;
    END
END AO21X1
MACRO AO21X2
    CLASS CORE ;
    FOREIGN AO21X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.65 4.90 0.75 9.60 ;
        RECT  0.25 5.40 0.75 9.60 ;
        RECT  0.25 9.10 1.80 9.60 ;
        RECT  0.65 4.90 1.15 6.30 ;
        RECT  0.25 5.40 1.15 6.30 ;
        RECT  1.10 9.10 1.80 9.80 ;
        RECT  0.65 4.90 2.55 5.40 ;
        RECT  2.05 2.75 2.55 5.40 ;
        RECT  2.05 2.75 2.75 3.45 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 3.95 5.35 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  5.45 5.40 6.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.55 7.30 2.75 7.80 ;
        RECT  1.55 7.10 2.25 7.80 ;
        RECT  2.25 7.30 2.75 11.00 ;
        RECT  5.90 7.75 6.60 11.00 ;
        RECT  0.00 11.00 8.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 4.45 ;
        RECT  3.40 2.00 4.10 3.45 ;
        RECT  7.25 2.00 7.95 4.50 ;
        RECT  0.00 0.00 8.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.40 5.85 3.70 6.60 ;
        RECT  3.20 5.85 3.70 10.55 ;
        RECT  3.20 7.20 3.90 10.55 ;
        RECT  4.45 4.00 4.95 6.35 ;
        RECT  4.90 2.70 4.95 6.35 ;
        RECT  2.40 5.85 4.95 6.35 ;
        RECT  4.55 6.80 5.25 10.55 ;
        RECT  4.90 2.70 5.60 4.50 ;
        RECT  4.45 4.00 5.60 4.50 ;
        RECT  4.55 6.80 7.95 7.30 ;
        RECT  7.25 6.80 7.95 10.55 ;
    END
END AO21X2
MACRO AO21X4
    CLASS CORE ;
    FOREIGN AO21X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  3.35 4.45 3.85 10.55 ;
        RECT  3.15 7.20 3.85 10.55 ;
        RECT  3.05 8.00 3.95 8.90 ;
        RECT  4.70 2.45 5.20 4.95 ;
        RECT  3.35 4.45 5.20 4.95 ;
        RECT  4.70 2.45 5.40 4.05 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  7.00 5.40 8.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  8.60 5.35 9.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.45 2.50 11.00 ;
        RECT  4.50 7.45 5.20 11.00 ;
        RECT  8.70 7.75 9.40 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 2.00 2.15 3.95 ;
        RECT  3.35 2.00 4.05 4.00 ;
        RECT  6.05 2.00 6.75 4.00 ;
        RECT  10.05 2.00 10.75 4.00 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.30 6.15 5.00 6.85 ;
        RECT  4.30 6.35 6.50 6.85 ;
        RECT  6.00 4.45 6.50 10.55 ;
        RECT  6.00 7.20 6.70 10.55 ;
        RECT  7.35 6.80 8.05 10.55 ;
        RECT  7.70 2.45 8.20 4.95 ;
        RECT  6.00 4.45 8.20 4.95 ;
        RECT  7.70 2.45 8.40 4.05 ;
        RECT  7.35 6.80 10.75 7.30 ;
        RECT  10.05 6.80 10.75 10.55 ;
    END
END AO21X4
MACRO AO221X1
    CLASS CORE ;
    FOREIGN AO221X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.30 3.00 11.10 3.70 ;
        RECT  10.60 3.00 11.10 9.40 ;
        RECT  10.40 7.70 11.10 9.40 ;
        RECT  10.40 8.00 12.35 8.90 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.35 8.15 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  5.50 4.10 6.75 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 3.95 5.00 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  1.65 4.10 2.55 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.50 7.55 4.20 11.00 ;
        RECT  9.05 7.70 9.75 11.00 ;
        RECT  9.05 10.35 12.15 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.25 2.00 1.95 3.65 ;
        RECT  5.95 2.00 6.65 2.70 ;
        RECT  8.95 2.00 9.65 3.70 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.00 5.55 1.50 10.55 ;
        RECT  0.80 8.15 1.50 10.55 ;
        RECT  2.15 6.55 2.85 10.55 ;
        RECT  3.60 2.55 4.30 3.65 ;
        RECT  2.15 6.55 5.55 7.05 ;
        RECT  4.85 6.55 5.55 10.55 ;
        RECT  1.00 5.55 6.70 6.05 ;
        RECT  6.20 5.55 6.70 10.55 ;
        RECT  6.20 6.75 6.90 10.55 ;
        RECT  3.60 3.15 8.15 3.65 ;
        RECT  7.45 3.00 8.15 3.75 ;
        RECT  7.65 3.00 8.15 4.85 ;
        RECT  7.55 6.75 8.25 10.55 ;
        RECT  7.65 4.35 10.15 4.85 ;
        RECT  8.65 4.35 9.15 7.25 ;
        RECT  7.55 6.75 9.15 7.25 ;
        RECT  8.65 4.35 10.15 5.05 ;
    END
END AO221X1
MACRO AO221X2
    CLASS CORE ;
    FOREIGN AO221X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.30 2.50 11.10 3.20 ;
        RECT  10.60 2.50 11.10 10.50 ;
        RECT  10.40 7.10 11.10 10.50 ;
        RECT  10.40 8.00 12.35 8.90 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.35 8.15 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  5.50 4.10 6.75 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 3.95 5.00 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  1.65 4.10 2.55 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.50 7.55 4.20 11.00 ;
        RECT  9.05 7.70 9.75 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.25 2.00 1.95 3.65 ;
        RECT  5.95 2.00 6.65 2.70 ;
        RECT  8.95 2.00 9.65 3.70 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.00 5.55 1.50 10.55 ;
        RECT  0.80 8.15 1.50 10.55 ;
        RECT  2.15 6.55 2.85 10.55 ;
        RECT  3.60 2.55 4.30 3.65 ;
        RECT  2.15 6.55 5.55 7.05 ;
        RECT  4.85 6.55 5.55 10.55 ;
        RECT  1.00 5.55 6.70 6.05 ;
        RECT  6.20 5.55 6.70 10.55 ;
        RECT  6.20 6.75 6.90 10.55 ;
        RECT  3.60 3.15 8.15 3.65 ;
        RECT  7.45 3.00 8.15 3.75 ;
        RECT  7.65 3.00 8.15 4.85 ;
        RECT  7.55 6.75 8.25 10.55 ;
        RECT  7.65 4.35 10.15 4.85 ;
        RECT  8.65 4.35 9.15 7.25 ;
        RECT  7.55 6.75 9.15 7.25 ;
        RECT  8.65 4.35 10.15 5.05 ;
    END
END AO221X2
MACRO AO221X4
    CLASS CORE ;
    FOREIGN AO221X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.40 5.60 10.90 10.50 ;
        RECT  10.40 7.10 11.10 10.50 ;
        RECT  11.50 2.45 12.20 4.05 ;
        RECT  11.70 2.45 12.20 6.10 ;
        RECT  10.40 5.60 12.20 6.10 ;
        RECT  11.45 2.80 12.35 3.70 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.35 8.15 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  5.50 4.10 6.75 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 3.95 5.00 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  1.65 4.10 2.55 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.50 7.45 4.20 11.00 ;
        RECT  9.05 7.70 9.75 11.00 ;
        RECT  11.75 7.70 12.45 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.25 2.00 1.95 3.65 ;
        RECT  5.95 2.00 6.65 2.70 ;
        RECT  10.15 2.00 10.85 3.95 ;
        RECT  12.85 2.00 13.55 3.95 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.00 5.55 1.50 10.55 ;
        RECT  0.80 8.15 1.50 10.55 ;
        RECT  2.15 6.50 2.85 10.55 ;
        RECT  3.60 2.55 4.30 3.65 ;
        RECT  2.15 6.50 5.55 7.00 ;
        RECT  4.85 6.50 5.55 10.55 ;
        RECT  1.00 5.55 6.70 6.05 ;
        RECT  6.20 5.55 6.70 10.55 ;
        RECT  6.20 6.75 6.90 10.55 ;
        RECT  3.60 3.15 8.15 3.65 ;
        RECT  7.45 3.00 8.15 3.75 ;
        RECT  7.65 3.00 8.15 4.90 ;
        RECT  7.55 6.75 8.25 10.55 ;
        RECT  8.65 4.40 9.15 7.25 ;
        RECT  7.55 6.75 9.15 7.25 ;
        RECT  7.65 4.40 11.20 4.90 ;
        RECT  10.50 4.40 11.20 5.10 ;
    END
END AO221X4
MACRO AO222X1
    CLASS CORE ;
    FOREIGN AO222X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.25 3.00 12.15 3.70 ;
        RECT  11.65 3.00 12.15 9.05 ;
        RECT  11.40 7.35 12.15 9.05 ;
        RECT  11.40 8.00 12.35 9.05 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.55 5.00 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  5.85 4.10 6.90 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  4.45 4.10 5.35 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 3.95 5.00 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  1.65 4.10 2.55 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.15 7.75 3.85 11.00 ;
        RECT  10.05 7.35 10.75 11.00 ;
        RECT  10.05 10.10 12.15 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.05 2.00 1.75 3.10 ;
        RECT  5.90 2.00 6.60 2.70 ;
        RECT  9.90 2.00 10.60 3.70 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.65 5.80 1.15 10.10 ;
        RECT  0.45 7.30 1.15 10.10 ;
        RECT  1.80 6.75 2.50 10.10 ;
        RECT  3.40 2.45 4.10 3.65 ;
        RECT  1.80 6.75 5.20 7.25 ;
        RECT  4.50 6.75 5.20 10.10 ;
        RECT  0.65 5.80 6.35 6.30 ;
        RECT  5.85 5.80 6.35 10.55 ;
        RECT  5.85 7.30 6.55 10.55 ;
        RECT  7.40 3.15 7.90 9.60 ;
        RECT  7.20 7.70 7.90 9.60 ;
        RECT  8.40 2.45 9.10 3.65 ;
        RECT  3.40 3.15 9.10 3.65 ;
        RECT  8.55 7.70 9.25 10.55 ;
        RECT  5.85 10.05 9.25 10.55 ;
        RECT  10.50 5.60 11.20 6.30 ;
        RECT  7.40 5.80 11.20 6.30 ;
    END
END AO222X1
MACRO AO222X2
    CLASS CORE ;
    FOREIGN AO222X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.40 2.45 12.15 4.05 ;
        RECT  11.65 2.45 12.10 10.50 ;
        RECT  11.40 7.10 12.10 10.50 ;
        RECT  11.65 2.45 12.15 8.90 ;
        RECT  11.40 7.10 12.15 8.90 ;
        RECT  11.40 8.00 12.35 8.90 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.55 5.00 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  5.85 4.10 6.90 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  4.45 4.10 5.35 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 3.95 5.00 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  1.65 4.10 2.55 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.15 7.75 3.85 11.00 ;
        RECT  10.05 7.10 10.75 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.05 2.00 1.75 3.10 ;
        RECT  5.90 2.00 6.60 2.70 ;
        RECT  9.90 2.00 10.60 3.70 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.65 5.80 1.15 10.10 ;
        RECT  0.45 7.30 1.15 10.10 ;
        RECT  1.80 6.75 2.50 10.10 ;
        RECT  3.40 2.45 4.10 3.65 ;
        RECT  1.80 6.75 5.20 7.25 ;
        RECT  4.50 6.75 5.20 10.10 ;
        RECT  0.65 5.80 6.35 6.30 ;
        RECT  5.85 5.80 6.35 10.55 ;
        RECT  5.85 7.30 6.55 10.55 ;
        RECT  7.40 3.15 7.90 9.60 ;
        RECT  7.20 7.70 7.90 9.60 ;
        RECT  8.40 2.45 9.10 3.65 ;
        RECT  3.40 3.15 9.10 3.65 ;
        RECT  8.55 7.70 9.25 10.55 ;
        RECT  5.85 10.05 9.25 10.55 ;
        RECT  10.50 5.60 11.20 6.30 ;
        RECT  7.40 5.80 11.20 6.30 ;
    END
END AO222X2
MACRO AO222X4
    CLASS CORE ;
    FOREIGN AO222X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.45 2.80 12.15 4.40 ;
        RECT  11.65 2.80 12.15 10.50 ;
        RECT  11.45 7.10 12.15 10.50 ;
        RECT  11.45 8.00 12.35 8.90 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.55 5.00 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  5.85 4.10 6.90 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  4.45 4.10 5.35 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 3.95 5.00 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  1.65 4.10 2.55 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.15 7.60 3.85 11.00 ;
        RECT  10.10 7.10 10.80 11.00 ;
        RECT  12.80 7.10 13.50 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.05 2.00 1.75 3.10 ;
        RECT  5.90 2.00 6.60 2.70 ;
        RECT  10.10 2.00 10.80 4.40 ;
        RECT  12.80 2.00 13.50 4.40 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.65 5.65 1.15 10.10 ;
        RECT  0.45 7.30 1.15 10.10 ;
        RECT  1.80 6.60 2.50 10.10 ;
        RECT  3.40 2.45 4.10 3.65 ;
        RECT  1.80 6.60 5.20 7.10 ;
        RECT  4.50 6.60 5.20 10.10 ;
        RECT  0.65 5.65 6.35 6.15 ;
        RECT  5.85 5.65 6.35 10.55 ;
        RECT  5.85 7.30 6.55 10.55 ;
        RECT  7.40 3.15 7.90 9.60 ;
        RECT  7.20 7.70 7.90 9.60 ;
        RECT  8.40 2.45 9.10 3.65 ;
        RECT  3.40 3.15 9.10 3.65 ;
        RECT  8.55 7.30 9.25 10.55 ;
        RECT  5.85 10.05 9.25 10.55 ;
        RECT  10.50 5.60 11.20 6.30 ;
        RECT  7.40 5.80 11.20 6.30 ;
    END
END AO222X4
MACRO AO22X1
    CLASS CORE ;
    FOREIGN AO22X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.25 3.15 0.75 10.40 ;
        RECT  0.25 9.30 1.15 10.40 ;
        RECT  1.20 2.95 1.90 3.65 ;
        RECT  0.25 3.15 1.90 3.65 ;
        RECT  0.25 9.70 3.45 10.40 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.20 5.40 5.35 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.20 5.40 8.15 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.55 4.10 6.75 4.80 ;
        RECT  5.85 4.10 6.75 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  5.90 7.80 6.60 11.00 ;
        RECT  4.40 10.10 7.95 11.00 ;
        RECT  0.00 11.00 8.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.55 2.00 3.25 3.65 ;
        RECT  7.25 2.00 7.95 3.65 ;
        RECT  0.00 0.00 8.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.65 4.10 2.35 4.80 ;
        RECT  1.85 7.20 2.55 9.25 ;
        RECT  3.20 4.30 3.70 8.30 ;
        RECT  3.20 7.60 3.90 8.30 ;
        RECT  3.80 3.15 4.30 4.80 ;
        RECT  1.65 4.30 4.30 4.80 ;
        RECT  4.55 6.85 5.25 9.25 ;
        RECT  1.85 8.75 5.25 9.25 ;
        RECT  4.90 2.95 5.60 3.65 ;
        RECT  3.80 3.15 5.60 3.65 ;
        RECT  4.55 6.85 7.95 7.35 ;
        RECT  7.25 6.85 7.95 8.90 ;
    END
END AO22X1
MACRO AO22X2
    CLASS CORE ;
    FOREIGN AO22X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.25 3.15 0.75 10.40 ;
        RECT  0.25 9.30 1.15 10.40 ;
        RECT  1.05 2.95 1.75 3.65 ;
        RECT  0.25 3.15 1.75 3.65 ;
        RECT  0.25 9.70 4.30 10.40 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.20 5.40 5.35 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.20 5.40 8.15 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.55 4.10 6.75 4.80 ;
        RECT  5.85 4.10 6.75 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  5.90 7.80 6.60 11.00 ;
        RECT  5.60 10.10 7.95 11.00 ;
        RECT  0.00 11.00 8.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.40 2.00 3.10 3.65 ;
        RECT  7.25 2.00 7.95 3.65 ;
        RECT  0.00 0.00 8.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.65 4.10 2.35 4.80 ;
        RECT  1.85 7.20 2.55 9.25 ;
        RECT  3.20 4.30 3.70 8.30 ;
        RECT  3.20 7.60 3.90 8.30 ;
        RECT  3.80 3.15 4.30 4.80 ;
        RECT  1.65 4.30 4.30 4.80 ;
        RECT  4.55 6.85 5.25 9.25 ;
        RECT  1.85 8.75 5.25 9.25 ;
        RECT  4.90 2.95 5.60 3.65 ;
        RECT  3.80 3.15 5.60 3.65 ;
        RECT  4.55 6.85 7.95 7.35 ;
        RECT  7.25 6.85 7.95 8.90 ;
    END
END AO22X2
MACRO AO22X4
    CLASS CORE ;
    FOREIGN AO22X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.65 9.30 2.55 10.20 ;
        RECT  2.05 4.80 2.55 10.55 ;
        RECT  1.80 7.15 2.55 10.55 ;
        RECT  3.70 2.65 4.40 5.30 ;
        RECT  2.05 4.80 4.40 5.30 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.35 7.60 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.20 5.40 8.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  10.00 5.40 10.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.40 9.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.35 1.15 11.00 ;
        RECT  3.15 7.35 3.85 11.00 ;
        RECT  8.70 8.10 9.40 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 2.00 1.20 4.40 ;
        RECT  2.35 2.00 3.05 4.35 ;
        RECT  5.05 2.00 5.75 4.35 ;
        RECT  9.90 2.00 10.60 4.35 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.25 5.75 3.95 6.50 ;
        RECT  4.65 8.05 5.35 10.45 ;
        RECT  3.25 5.75 6.70 6.25 ;
        RECT  6.20 3.85 6.70 9.50 ;
        RECT  6.00 7.90 6.70 9.50 ;
        RECT  7.35 7.15 8.05 10.45 ;
        RECT  4.65 9.95 8.05 10.45 ;
        RECT  7.55 3.65 8.25 4.35 ;
        RECT  6.20 3.85 8.25 4.35 ;
        RECT  7.35 7.15 10.75 7.65 ;
        RECT  10.05 7.15 10.75 9.55 ;
    END
END AO22X4
MACRO AO311X1
    CLASS CORE ;
    FOREIGN AO311X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.50 3.00 1.00 10.20 ;
        RECT  0.50 7.15 1.20 10.20 ;
        RECT  0.25 9.30 1.20 10.20 ;
        RECT  0.50 3.00 2.05 3.70 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.55 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  7.25 4.10 8.15 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  5.85 4.10 6.75 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  4.30 5.35 5.35 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.35 3.30 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.00 7.10 2.70 11.00 ;
        RECT  4.70 7.70 5.40 11.00 ;
        RECT  9.95 9.55 10.65 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.85 2.00 3.55 3.70 ;
        RECT  7.70 2.00 8.40 2.70 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.45 4.15 2.15 4.85 ;
        RECT  3.35 6.75 4.05 10.55 ;
        RECT  4.15 3.15 4.65 4.65 ;
        RECT  1.45 4.15 4.65 4.65 ;
        RECT  3.35 6.75 6.75 7.25 ;
        RECT  6.05 6.40 6.75 10.55 ;
        RECT  6.20 2.45 6.90 3.65 ;
        RECT  8.40 6.40 9.10 10.20 ;
        RECT  9.20 2.45 9.90 3.65 ;
        RECT  4.15 3.15 10.50 3.65 ;
        RECT  10.00 3.15 10.50 6.90 ;
        RECT  8.40 6.40 10.50 6.90 ;
    END
END AO311X1
MACRO AO311X2
    CLASS CORE ;
    FOREIGN AO311X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.50 3.00 1.00 10.55 ;
        RECT  0.50 7.10 1.20 10.55 ;
        RECT  0.25 9.30 1.20 10.55 ;
        RECT  0.50 3.00 2.05 3.70 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.55 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  7.25 4.10 8.15 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  5.85 4.10 6.75 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  4.30 5.35 5.35 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.35 3.30 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.00 7.10 2.70 11.00 ;
        RECT  4.70 7.70 5.40 11.00 ;
        RECT  9.95 9.55 10.65 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.85 2.00 3.55 3.70 ;
        RECT  7.70 2.00 8.40 2.70 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.45 4.15 2.15 4.85 ;
        RECT  3.35 6.75 4.05 10.55 ;
        RECT  4.15 3.15 4.65 4.65 ;
        RECT  1.45 4.15 4.65 4.65 ;
        RECT  3.35 6.75 6.75 7.25 ;
        RECT  6.05 6.40 6.75 10.55 ;
        RECT  6.20 2.45 6.90 3.65 ;
        RECT  8.40 6.40 9.10 10.20 ;
        RECT  9.20 2.45 9.90 3.65 ;
        RECT  4.15 3.15 10.50 3.65 ;
        RECT  10.00 3.15 10.50 6.90 ;
        RECT  8.40 6.40 10.50 6.90 ;
    END
END AO311X2
MACRO AO311X4
    CLASS CORE ;
    FOREIGN AO311X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.65 2.95 2.60 3.70 ;
        RECT  2.10 2.80 2.55 10.55 ;
        RECT  1.65 2.80 2.55 3.70 ;
        RECT  2.10 2.95 2.60 10.55 ;
        RECT  1.90 7.10 2.60 10.55 ;
        RECT  1.65 2.95 3.85 3.65 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  10.05 4.10 10.95 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.55 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  7.25 4.10 8.15 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  5.70 5.35 6.75 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.35 5.00 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.55 7.10 1.25 11.00 ;
        RECT  3.40 7.10 4.10 11.00 ;
        RECT  6.10 7.70 6.80 11.00 ;
        RECT  11.35 9.55 12.05 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 2.00 1.20 3.80 ;
        RECT  3.15 2.00 5.20 2.30 ;
        RECT  4.50 2.00 5.20 3.65 ;
        RECT  9.35 2.00 10.05 2.70 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.60 4.10 4.30 4.80 ;
        RECT  4.75 6.75 5.45 10.55 ;
        RECT  5.75 3.15 6.25 4.65 ;
        RECT  3.60 4.10 6.25 4.65 ;
        RECT  4.75 6.75 8.15 7.25 ;
        RECT  7.45 6.40 8.15 10.55 ;
        RECT  7.85 2.45 8.55 3.65 ;
        RECT  9.80 6.40 10.50 10.20 ;
        RECT  5.75 3.15 11.90 3.65 ;
        RECT  11.40 2.45 11.55 6.90 ;
        RECT  10.85 2.45 11.55 3.65 ;
        RECT  11.40 3.15 11.90 6.90 ;
        RECT  9.80 6.40 11.90 6.90 ;
    END
END AO311X4
MACRO AO31X1
    CLASS CORE ;
    FOREIGN AO31X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.40 3.75 0.90 10.25 ;
        RECT  0.40 3.75 1.15 4.45 ;
        RECT  0.40 7.30 1.15 10.25 ;
        RECT  0.25 9.25 1.25 10.25 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  5.80 5.40 6.75 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  4.05 5.40 5.35 6.35 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  2.05 6.15 2.55 7.60 ;
        RECT  1.65 6.70 2.55 7.60 ;
        RECT  2.05 6.15 3.10 6.85 ;
        RECT  1.65 6.70 3.10 6.85 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.95 8.05 2.65 11.00 ;
        RECT  4.65 8.25 5.35 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.95 2.00 2.65 4.50 ;
        RECT  6.80 2.00 7.50 3.60 ;
        RECT  8.65 2.00 9.35 3.80 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.35 4.95 2.05 5.65 ;
        RECT  3.10 4.25 3.60 5.45 ;
        RECT  1.35 4.95 3.60 5.45 ;
        RECT  3.30 7.30 4.00 10.55 ;
        RECT  3.30 7.30 6.70 7.80 ;
        RECT  5.30 2.45 6.00 4.75 ;
        RECT  6.00 7.30 6.70 10.55 ;
        RECT  7.35 7.30 8.05 10.55 ;
        RECT  3.10 4.25 9.10 4.75 ;
        RECT  8.60 4.25 9.10 7.80 ;
        RECT  7.35 7.30 9.10 7.80 ;
    END
END AO31X1
MACRO AO31X2
    CLASS CORE ;
    FOREIGN AO31X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.40 2.75 0.90 10.20 ;
        RECT  0.40 2.75 1.15 4.45 ;
        RECT  0.40 7.30 1.15 10.20 ;
        RECT  0.25 9.25 1.15 10.20 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  5.80 5.35 6.75 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  4.05 5.40 5.35 6.35 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  2.05 6.15 2.55 7.60 ;
        RECT  1.65 6.70 2.55 7.60 ;
        RECT  2.05 6.15 3.10 6.85 ;
        RECT  1.65 6.70 3.10 6.85 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.05 2.50 11.00 ;
        RECT  4.50 8.25 5.20 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.95 2.00 2.65 4.50 ;
        RECT  6.80 2.00 7.50 3.60 ;
        RECT  8.65 2.00 9.35 3.80 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.35 4.95 2.05 5.65 ;
        RECT  3.10 4.25 3.60 5.45 ;
        RECT  1.35 4.95 3.60 5.45 ;
        RECT  3.15 7.30 3.85 10.55 ;
        RECT  3.15 7.30 6.55 7.80 ;
        RECT  5.30 2.45 6.00 4.75 ;
        RECT  5.85 7.30 6.55 10.55 ;
        RECT  7.20 7.30 7.90 10.55 ;
        RECT  3.10 4.25 9.10 4.75 ;
        RECT  8.60 4.25 9.10 7.80 ;
        RECT  7.20 7.30 9.10 7.80 ;
    END
END AO31X2
MACRO AO31X4
    CLASS CORE ;
    FOREIGN AO31X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.45 2.30 10.55 ;
        RECT  1.80 2.45 2.50 4.05 ;
        RECT  1.80 7.15 2.50 10.55 ;
        RECT  1.65 9.30 2.55 10.55 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.55 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  7.20 5.25 8.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  5.60 5.40 6.75 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.45 6.05 3.95 7.60 ;
        RECT  3.05 6.70 3.95 7.60 ;
        RECT  3.45 6.05 4.20 6.75 ;
        RECT  3.05 6.70 4.20 6.75 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.20 1.15 11.00 ;
        RECT  3.15 8.05 3.85 11.00 ;
        RECT  5.85 8.65 6.55 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 4.05 ;
        RECT  3.15 2.00 3.85 3.90 ;
        RECT  8.00 2.00 8.70 3.65 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.75 4.45 3.45 5.15 ;
        RECT  2.75 4.65 5.15 5.15 ;
        RECT  4.65 4.15 5.15 7.25 ;
        RECT  4.50 7.70 5.20 10.55 ;
        RECT  4.65 4.15 7.20 4.65 ;
        RECT  4.50 7.70 7.90 8.20 ;
        RECT  6.50 2.45 7.20 4.65 ;
        RECT  7.20 7.70 7.90 10.55 ;
        RECT  4.65 6.75 9.25 7.25 ;
        RECT  8.55 6.75 9.25 10.55 ;
    END
END AO31X4
MACRO AO321X1
    CLASS CORE ;
    FOREIGN AO321X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.45 3.20 0.95 10.20 ;
        RECT  0.45 7.15 1.15 10.20 ;
        RECT  0.25 9.30 1.15 10.20 ;
        RECT  1.70 3.00 2.40 3.70 ;
        RECT  0.45 3.20 2.40 3.70 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  11.45 4.10 12.35 5.00 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  7.25 4.10 8.15 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.55 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  5.85 4.10 6.75 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  4.30 5.10 5.35 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.35 3.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.95 7.10 2.65 11.00 ;
        RECT  4.65 7.70 5.35 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.25 2.00 3.95 3.70 ;
        RECT  8.95 2.00 10.55 2.70 ;
        RECT  12.85 2.00 13.55 3.80 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.40 4.15 2.10 4.85 ;
        RECT  3.30 6.75 4.00 10.55 ;
        RECT  4.55 3.15 5.05 4.65 ;
        RECT  1.40 4.15 5.05 4.65 ;
        RECT  3.30 6.75 6.70 7.25 ;
        RECT  6.00 6.40 6.70 10.55 ;
        RECT  6.60 2.55 7.30 3.65 ;
        RECT  7.35 6.40 8.05 9.60 ;
        RECT  8.70 7.35 9.40 10.55 ;
        RECT  6.00 10.05 9.40 10.55 ;
        RECT  7.35 6.40 10.90 6.90 ;
        RECT  10.20 3.15 10.70 5.95 ;
        RECT  10.20 6.40 10.90 10.55 ;
        RECT  10.20 5.45 12.25 5.95 ;
        RECT  11.35 2.45 12.05 3.65 ;
        RECT  4.55 3.15 12.05 3.65 ;
        RECT  11.55 5.45 12.25 10.20 ;
    END
END AO321X1
MACRO AO321X2
    CLASS CORE ;
    FOREIGN AO321X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.80 0.95 10.50 ;
        RECT  0.45 7.10 1.15 10.50 ;
        RECT  0.25 9.30 1.15 10.50 ;
        RECT  1.70 2.60 2.40 3.30 ;
        RECT  0.45 2.80 2.40 3.30 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  11.45 4.10 12.35 5.00 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  7.25 4.10 8.15 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.55 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  5.85 4.10 6.75 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  4.30 5.10 5.35 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.35 3.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.95 7.10 2.65 11.00 ;
        RECT  4.65 7.70 5.35 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.25 2.00 3.95 3.70 ;
        RECT  8.95 2.00 10.55 2.70 ;
        RECT  12.85 2.00 13.55 3.80 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.40 4.15 2.10 4.85 ;
        RECT  3.30 6.75 4.00 10.55 ;
        RECT  4.55 3.15 5.05 4.65 ;
        RECT  1.40 4.15 5.05 4.65 ;
        RECT  3.30 6.75 6.70 7.25 ;
        RECT  6.00 6.40 6.70 10.55 ;
        RECT  6.60 2.55 7.30 3.65 ;
        RECT  7.35 6.40 8.05 9.60 ;
        RECT  8.70 7.35 9.40 10.55 ;
        RECT  6.00 10.05 9.40 10.55 ;
        RECT  7.35 6.40 10.90 6.90 ;
        RECT  10.20 3.15 10.70 5.95 ;
        RECT  10.20 6.40 10.90 10.55 ;
        RECT  10.20 5.45 12.25 5.95 ;
        RECT  11.35 2.45 12.05 3.65 ;
        RECT  4.55 3.15 12.05 3.65 ;
        RECT  11.55 5.45 12.25 10.20 ;
    END
END AO321X2
MACRO AO321X4
    CLASS CORE ;
    FOREIGN AO321X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.80 2.30 10.50 ;
        RECT  1.80 7.10 2.50 10.50 ;
        RECT  1.65 2.80 2.55 3.70 ;
        RECT  1.65 3.00 3.65 3.70 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  12.85 4.10 13.75 5.00 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.55 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  10.05 4.10 10.95 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  7.25 4.10 8.15 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  5.50 5.10 6.75 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.35 4.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.10 1.15 11.00 ;
        RECT  3.15 7.10 3.85 11.00 ;
        RECT  5.85 7.70 6.55 11.00 ;
        RECT  14.25 9.55 14.95 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 2.00 1.20 3.60 ;
        RECT  0.50 2.00 2.65 2.35 ;
        RECT  4.45 2.00 5.15 3.70 ;
        RECT  10.35 2.00 11.95 2.70 ;
        RECT  14.25 2.00 14.95 3.80 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.80 4.15 3.50 4.85 ;
        RECT  4.50 6.75 5.20 10.55 ;
        RECT  5.95 3.15 6.45 4.65 ;
        RECT  2.80 4.15 6.45 4.65 ;
        RECT  4.50 6.75 7.90 7.25 ;
        RECT  7.20 6.40 7.90 10.55 ;
        RECT  7.80 2.55 8.50 3.65 ;
        RECT  8.55 6.40 9.25 9.60 ;
        RECT  9.90 7.35 10.60 10.55 ;
        RECT  7.20 10.05 10.60 10.55 ;
        RECT  8.55 6.40 12.10 6.90 ;
        RECT  11.60 3.15 12.10 5.95 ;
        RECT  11.40 6.40 12.10 10.55 ;
        RECT  11.60 5.45 13.45 5.95 ;
        RECT  12.75 2.45 13.45 3.65 ;
        RECT  5.95 3.15 13.45 3.65 ;
        RECT  12.75 5.45 13.45 10.55 ;
    END
END AO321X4
MACRO AO322X1
    CLASS CORE ;
    FOREIGN AO322X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.55 0.95 10.20 ;
        RECT  0.45 2.55 1.15 3.25 ;
        RECT  0.45 7.75 1.15 10.20 ;
        RECT  0.25 9.30 1.15 10.20 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  10.05 4.10 10.95 5.00 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.40 9.55 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  7.25 4.10 8.15 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  4.45 4.10 5.35 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 4.20 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.75 2.50 11.00 ;
        RECT  4.50 7.70 5.20 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 3.25 ;
        RECT  7.65 2.00 8.35 2.70 ;
        RECT  12.75 2.00 13.55 3.80 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.40 3.75 2.10 4.45 ;
        RECT  3.10 3.15 3.60 4.25 ;
        RECT  1.40 3.75 3.60 4.25 ;
        RECT  3.15 6.75 3.85 10.50 ;
        RECT  3.15 6.75 6.55 7.25 ;
        RECT  5.15 2.50 5.85 3.65 ;
        RECT  5.85 6.75 6.55 10.55 ;
        RECT  7.20 6.75 7.90 9.60 ;
        RECT  8.55 7.70 9.25 10.55 ;
        RECT  5.85 10.05 9.25 10.55 ;
        RECT  7.20 6.75 10.75 7.25 ;
        RECT  10.05 6.75 10.75 10.55 ;
        RECT  10.15 2.55 10.85 3.65 ;
        RECT  3.10 3.15 11.90 3.65 ;
        RECT  11.40 3.15 11.90 9.60 ;
        RECT  11.40 7.70 12.10 9.60 ;
        RECT  12.75 7.70 13.45 10.55 ;
        RECT  10.05 10.05 13.45 10.55 ;
    END
END AO322X1
MACRO AO322X2
    CLASS CORE ;
    FOREIGN AO322X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.55 0.95 10.45 ;
        RECT  0.45 2.55 1.15 3.25 ;
        RECT  0.45 7.55 1.15 10.45 ;
        RECT  0.25 9.30 1.15 10.45 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  10.05 4.10 10.95 5.00 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.40 9.55 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  7.25 4.10 8.15 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  4.45 4.10 5.35 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 4.20 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.35 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.75 2.50 11.00 ;
        RECT  4.50 7.70 5.20 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 3.05 ;
        RECT  7.65 2.00 8.35 2.70 ;
        RECT  12.75 2.00 13.55 3.80 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.40 4.10 2.10 4.80 ;
        RECT  3.10 3.15 3.60 4.60 ;
        RECT  1.40 4.10 3.60 4.60 ;
        RECT  3.15 6.75 3.85 10.50 ;
        RECT  3.15 6.75 6.55 7.25 ;
        RECT  5.15 2.50 5.85 3.65 ;
        RECT  5.85 6.75 6.55 10.55 ;
        RECT  7.20 6.75 7.90 9.60 ;
        RECT  8.55 7.70 9.25 10.55 ;
        RECT  5.85 10.05 9.25 10.55 ;
        RECT  7.20 6.75 10.75 7.25 ;
        RECT  10.05 6.75 10.75 10.55 ;
        RECT  10.15 2.55 10.85 3.65 ;
        RECT  3.10 3.15 11.90 3.65 ;
        RECT  11.40 3.15 11.90 9.60 ;
        RECT  11.40 7.70 12.10 9.60 ;
        RECT  12.75 7.70 13.45 10.55 ;
        RECT  10.05 10.05 13.45 10.55 ;
    END
END AO322X2
MACRO AO322X4
    CLASS CORE ;
    FOREIGN AO322X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.45 2.30 10.55 ;
        RECT  1.80 2.45 2.50 4.05 ;
        RECT  1.80 7.75 2.55 10.55 ;
        RECT  1.65 9.30 2.55 10.55 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  11.45 4.10 12.35 5.00 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.55 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  5.85 4.10 6.75 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        RECT  4.45 5.50 5.80 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 4.20 7.60 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 8.10 1.15 11.00 ;
        RECT  3.15 8.10 3.85 11.00 ;
        RECT  6.00 7.75 6.70 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.95 ;
        RECT  3.15 2.00 3.85 3.95 ;
        RECT  9.15 2.00 9.85 2.70 ;
        RECT  13.20 2.00 14.80 2.20 ;
        RECT  14.10 2.00 14.80 3.30 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.80 4.40 3.50 5.10 ;
        RECT  4.50 3.15 5.00 4.90 ;
        RECT  2.80 4.40 5.00 4.90 ;
        RECT  4.65 6.75 5.35 10.50 ;
        RECT  4.65 6.75 8.05 7.25 ;
        RECT  6.65 2.50 7.35 3.65 ;
        RECT  7.35 6.75 8.05 10.55 ;
        RECT  8.70 6.75 9.40 9.60 ;
        RECT  10.05 7.75 10.75 10.55 ;
        RECT  7.35 10.05 10.75 10.55 ;
        RECT  8.70 6.75 12.25 7.25 ;
        RECT  11.55 6.75 12.25 10.55 ;
        RECT  11.65 2.55 12.35 3.65 ;
        RECT  4.50 3.15 13.40 3.65 ;
        RECT  12.90 3.15 13.40 9.60 ;
        RECT  12.90 7.10 13.60 9.60 ;
        RECT  14.25 7.10 14.95 10.55 ;
        RECT  11.55 10.05 14.95 10.55 ;
    END
END AO322X4
MACRO AO32X1
    CLASS CORE ;
    FOREIGN AO32X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.25 3.40 0.75 10.20 ;
        RECT  0.25 3.40 1.15 4.10 ;
        RECT  0.25 8.05 1.15 10.20 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.55 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 4.00 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.55 7.60 ;
        RECT  1.65 6.85 2.85 7.60 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.05 2.50 11.00 ;
        RECT  4.50 8.05 5.20 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.95 2.00 2.65 3.90 ;
        RECT  7.65 2.00 8.35 3.65 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.45 4.45 1.95 5.25 ;
        RECT  1.25 4.55 1.95 5.25 ;
        RECT  3.35 7.05 3.85 9.75 ;
        RECT  3.15 8.05 3.85 9.75 ;
        RECT  3.35 7.05 6.55 7.55 ;
        RECT  5.30 2.90 6.00 4.95 ;
        RECT  5.85 7.05 6.55 10.55 ;
        RECT  1.45 4.45 7.70 4.95 ;
        RECT  1.25 4.55 7.70 4.95 ;
        RECT  7.20 4.45 7.70 9.60 ;
        RECT  7.20 8.00 7.90 9.60 ;
        RECT  8.55 8.05 9.25 10.55 ;
        RECT  5.85 10.05 9.25 10.55 ;
    END
END AO32X1
MACRO AO32X2
    CLASS CORE ;
    FOREIGN AO32X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.25 2.50 0.75 10.50 ;
        RECT  0.25 2.50 1.15 4.10 ;
        RECT  0.25 8.00 1.15 10.50 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.55 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 4.00 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.55 7.60 ;
        RECT  1.65 6.85 2.85 7.60 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.05 2.50 11.00 ;
        RECT  4.50 8.05 5.20 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.00 ;
        RECT  7.65 2.00 8.35 3.65 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.45 4.45 1.95 5.25 ;
        RECT  1.25 4.55 1.95 5.25 ;
        RECT  3.35 7.05 3.85 9.75 ;
        RECT  3.15 8.05 3.85 9.75 ;
        RECT  3.35 7.05 6.55 7.55 ;
        RECT  5.30 2.90 6.00 4.95 ;
        RECT  5.85 7.05 6.55 10.55 ;
        RECT  1.45 4.45 7.70 4.95 ;
        RECT  1.25 4.55 7.70 4.95 ;
        RECT  7.20 4.45 7.70 9.60 ;
        RECT  7.20 8.00 7.90 9.60 ;
        RECT  8.55 8.05 9.25 10.55 ;
        RECT  5.85 10.05 9.25 10.55 ;
    END
END AO32X2
MACRO AO32X4
    CLASS CORE ;
    FOREIGN AO32X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.50 2.20 10.50 ;
        RECT  1.70 3.60 2.20 10.50 ;
        RECT  1.80 2.50 2.50 4.10 ;
        RECT  1.70 3.60 2.50 4.10 ;
        RECT  1.70 8.00 2.55 10.50 ;
        RECT  1.65 9.30 2.55 10.50 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  10.05 4.10 10.95 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.40 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        RECT  3.05 6.85 4.20 7.60 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 8.05 1.15 11.00 ;
        RECT  3.15 8.05 3.85 11.00 ;
        RECT  6.00 8.05 6.70 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 4.00 ;
        RECT  3.15 2.00 3.85 4.00 ;
        RECT  9.00 2.00 9.70 3.65 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.85 4.45 3.35 5.25 ;
        RECT  2.65 4.55 3.35 5.25 ;
        RECT  4.85 7.05 5.35 9.75 ;
        RECT  4.65 8.05 5.35 9.75 ;
        RECT  4.85 7.05 8.05 7.55 ;
        RECT  6.65 2.90 7.35 4.95 ;
        RECT  7.35 7.05 8.05 10.55 ;
        RECT  2.85 4.45 9.20 4.95 ;
        RECT  2.65 4.55 9.20 4.95 ;
        RECT  8.70 4.45 9.20 9.60 ;
        RECT  8.70 8.00 9.40 9.60 ;
        RECT  10.05 8.05 10.75 10.55 ;
        RECT  7.35 10.05 10.75 10.55 ;
    END
END AO32X4
MACRO AO331X1
    CLASS CORE ;
    FOREIGN AO331X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.40 2.80 13.75 3.60 ;
        RECT  12.15 2.80 12.65 9.00 ;
        RECT  11.95 7.30 12.65 9.00 ;
        RECT  12.15 2.80 13.75 3.70 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  1.65 4.10 2.55 5.00 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  5.85 4.10 6.75 5.00 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  4.45 4.10 5.35 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 3.95 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  7.20 4.10 8.15 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  8.50 5.30 9.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  10.00 5.30 10.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  7.75 7.70 8.45 11.00 ;
        RECT  10.45 6.85 11.15 11.00 ;
        RECT  11.95 10.10 13.55 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.90 2.00 3.60 2.70 ;
        RECT  9.90 2.00 10.60 3.55 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.65 8.10 1.70 8.60 ;
        RECT  1.00 3.15 1.15 10.55 ;
        RECT  0.65 3.15 1.15 8.60 ;
        RECT  1.00 8.10 1.70 10.55 ;
        RECT  1.40 2.90 2.10 3.65 ;
        RECT  2.35 5.45 3.05 10.55 ;
        RECT  3.70 6.40 4.40 10.55 ;
        RECT  2.35 5.45 5.75 5.95 ;
        RECT  5.05 5.45 5.75 9.60 ;
        RECT  6.40 2.45 7.10 3.65 ;
        RECT  6.40 6.75 7.10 10.55 ;
        RECT  3.70 10.05 7.10 10.55 ;
        RECT  0.65 3.15 9.30 3.65 ;
        RECT  6.40 6.75 9.80 7.25 ;
        RECT  8.80 3.15 9.30 4.55 ;
        RECT  9.10 6.75 9.80 10.55 ;
        RECT  8.80 4.05 11.65 4.55 ;
        RECT  10.95 4.05 11.65 4.75 ;
    END
END AO331X1
MACRO AO331X2
    CLASS CORE ;
    FOREIGN AO331X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.40 2.80 13.75 3.60 ;
        RECT  12.15 2.80 12.65 10.50 ;
        RECT  11.95 7.10 12.65 10.50 ;
        RECT  12.15 2.80 13.75 3.70 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  1.65 4.10 2.55 5.00 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  5.85 4.10 6.75 5.00 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  4.45 4.10 5.35 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 3.95 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  7.20 4.10 8.15 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  8.50 5.30 9.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  10.00 5.30 10.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  7.75 7.70 8.45 11.00 ;
        RECT  10.45 6.85 11.15 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.90 2.00 3.60 2.70 ;
        RECT  9.90 2.00 10.60 3.55 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.65 8.10 1.70 8.60 ;
        RECT  1.00 3.15 1.15 10.55 ;
        RECT  0.65 3.15 1.15 8.60 ;
        RECT  1.00 8.10 1.70 10.55 ;
        RECT  1.40 2.90 2.10 3.65 ;
        RECT  2.35 5.45 3.05 10.55 ;
        RECT  3.70 6.40 4.40 10.55 ;
        RECT  2.35 5.45 5.75 5.95 ;
        RECT  5.05 5.45 5.75 9.60 ;
        RECT  6.40 2.45 7.10 3.65 ;
        RECT  6.40 6.75 7.10 10.55 ;
        RECT  3.70 10.05 7.10 10.55 ;
        RECT  0.65 3.15 9.30 3.65 ;
        RECT  6.40 6.75 9.80 7.25 ;
        RECT  8.80 3.15 9.30 4.55 ;
        RECT  9.10 6.75 9.80 10.55 ;
        RECT  8.80 4.05 11.65 4.55 ;
        RECT  10.95 4.05 11.65 4.75 ;
    END
END AO331X2
MACRO AO331X4
    CLASS CORE ;
    FOREIGN AO331X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  12.15 2.90 12.65 10.55 ;
        RECT  11.95 7.10 12.65 10.55 ;
        RECT  11.25 2.90 13.40 3.60 ;
        RECT  12.15 5.40 13.75 6.30 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  1.65 4.10 2.55 5.00 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  5.85 4.10 6.75 5.00 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  4.45 4.10 5.35 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 3.95 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  7.20 4.10 8.15 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  8.50 5.30 9.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  10.00 5.30 10.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  7.75 7.70 8.45 11.00 ;
        RECT  10.45 7.10 11.15 11.00 ;
        RECT  13.30 7.10 14.00 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.90 2.00 3.60 2.70 ;
        RECT  9.90 2.00 10.60 3.55 ;
        RECT  9.90 2.00 12.40 2.25 ;
        RECT  14.25 2.00 14.95 3.80 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.65 8.10 1.70 8.60 ;
        RECT  1.00 3.15 1.15 10.55 ;
        RECT  0.65 3.15 1.15 8.60 ;
        RECT  1.00 8.10 1.70 10.55 ;
        RECT  1.40 2.90 2.10 3.65 ;
        RECT  2.35 5.45 3.05 10.55 ;
        RECT  3.70 6.40 4.40 10.55 ;
        RECT  2.35 5.45 5.75 5.95 ;
        RECT  5.05 5.45 5.75 9.60 ;
        RECT  6.40 2.45 7.10 3.65 ;
        RECT  6.40 6.75 7.10 10.55 ;
        RECT  3.70 10.05 7.10 10.55 ;
        RECT  0.65 3.15 9.30 3.65 ;
        RECT  6.40 6.75 9.80 7.25 ;
        RECT  8.80 3.15 9.30 4.55 ;
        RECT  9.10 6.75 9.80 10.55 ;
        RECT  8.80 4.05 11.50 4.55 ;
        RECT  10.80 4.05 11.50 4.75 ;
    END
END AO331X4
MACRO AO332X1
    CLASS CORE ;
    FOREIGN AO332X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.55 0.95 10.20 ;
        RECT  0.45 2.55 1.15 3.25 ;
        RECT  0.45 7.75 1.15 10.20 ;
        RECT  0.25 9.30 1.15 10.20 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  8.45 4.10 9.55 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  4.45 4.10 5.35 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 4.20 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.75 2.50 11.00 ;
        RECT  4.50 7.70 5.20 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 3.25 ;
        RECT  8.65 2.00 9.35 2.70 ;
        RECT  12.75 2.00 13.55 3.80 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.40 3.75 2.10 4.45 ;
        RECT  3.10 3.15 3.60 4.25 ;
        RECT  1.40 3.75 3.60 4.25 ;
        RECT  3.15 6.75 3.85 10.50 ;
        RECT  3.15 6.75 6.55 7.25 ;
        RECT  5.15 2.50 5.85 3.65 ;
        RECT  5.85 6.75 6.55 10.55 ;
        RECT  7.20 6.75 7.90 9.60 ;
        RECT  8.55 7.70 9.25 10.55 ;
        RECT  5.85 10.05 9.25 10.55 ;
        RECT  7.20 6.75 10.60 7.25 ;
        RECT  9.90 6.75 10.60 10.55 ;
        RECT  11.15 2.55 11.95 3.65 ;
        RECT  3.10 3.15 11.95 3.65 ;
        RECT  11.45 2.55 11.95 9.60 ;
        RECT  11.25 7.70 11.95 9.60 ;
        RECT  12.60 7.70 13.30 10.55 ;
        RECT  9.90 10.05 13.30 10.55 ;
    END
END AO332X1
MACRO AO332X2
    CLASS CORE ;
    FOREIGN AO332X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.55 0.95 10.20 ;
        RECT  0.45 2.55 1.15 3.25 ;
        RECT  0.45 7.30 1.15 10.20 ;
        RECT  0.25 9.30 1.15 10.20 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  8.45 4.10 9.55 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  4.45 4.10 5.35 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 4.20 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.70 2.50 11.00 ;
        RECT  4.50 7.70 5.20 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 3.25 ;
        RECT  8.65 2.00 9.35 2.70 ;
        RECT  12.75 2.00 13.55 3.80 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.40 3.75 2.10 4.45 ;
        RECT  3.10 3.15 3.60 4.25 ;
        RECT  1.40 3.75 3.60 4.25 ;
        RECT  3.15 6.75 3.85 10.50 ;
        RECT  3.15 6.75 6.55 7.25 ;
        RECT  5.15 2.50 5.85 3.65 ;
        RECT  5.85 6.75 6.55 10.55 ;
        RECT  7.20 6.75 7.90 9.60 ;
        RECT  8.55 7.70 9.25 10.55 ;
        RECT  5.85 10.05 9.25 10.55 ;
        RECT  7.20 6.75 10.60 7.25 ;
        RECT  9.90 6.75 10.60 10.55 ;
        RECT  11.15 2.55 11.95 3.65 ;
        RECT  3.10 3.15 11.95 3.65 ;
        RECT  11.45 2.55 11.95 9.60 ;
        RECT  11.25 7.70 11.95 9.60 ;
        RECT  12.60 7.70 13.30 10.55 ;
        RECT  9.90 10.05 13.30 10.55 ;
    END
END AO332X2
MACRO AO332X4
    CLASS CORE ;
    FOREIGN AO332X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.45 2.30 10.55 ;
        RECT  1.80 2.45 2.50 4.05 ;
        RECT  1.80 7.85 2.55 10.55 ;
        RECT  1.65 9.30 2.55 10.55 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.40 9.55 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  9.95 4.10 10.95 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  5.85 4.10 6.75 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        RECT  4.45 5.55 5.70 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        RECT  3.05 6.75 4.25 7.60 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 8.05 1.15 11.00 ;
        RECT  3.15 8.05 3.85 11.00 ;
        RECT  6.00 7.80 6.70 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.95 ;
        RECT  3.15 2.00 3.85 3.95 ;
        RECT  10.15 2.00 10.85 2.70 ;
        RECT  14.15 2.00 14.85 3.50 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.80 4.40 3.50 5.10 ;
        RECT  4.50 3.15 5.00 4.90 ;
        RECT  2.80 4.40 5.00 4.90 ;
        RECT  4.80 6.75 5.35 10.55 ;
        RECT  4.65 8.05 5.35 10.55 ;
        RECT  4.80 6.75 8.05 7.25 ;
        RECT  6.65 2.50 7.35 3.65 ;
        RECT  7.35 6.75 8.05 10.55 ;
        RECT  8.70 6.75 9.40 9.60 ;
        RECT  10.05 7.80 10.75 10.55 ;
        RECT  7.35 10.05 10.75 10.55 ;
        RECT  8.70 6.75 12.10 7.25 ;
        RECT  11.40 6.75 12.10 10.55 ;
        RECT  12.65 2.85 13.45 3.65 ;
        RECT  4.50 3.15 13.45 3.65 ;
        RECT  12.95 2.85 13.45 9.60 ;
        RECT  12.75 7.80 13.45 9.60 ;
        RECT  14.10 7.80 14.80 10.55 ;
        RECT  11.40 10.05 14.80 10.55 ;
    END
END AO332X4
MACRO AO333X1
    CLASS CORE ;
    FOREIGN AO333X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.95 0.95 10.20 ;
        RECT  0.45 2.95 1.15 3.65 ;
        RECT  0.45 7.75 1.15 10.20 ;
        RECT  0.25 9.30 1.15 10.20 ;
        END
    END Q
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  12.85 4.10 13.75 5.00 ;
        END
    END J
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  10.05 4.10 10.95 5.00 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.40 9.55 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 4.10 5.35 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        RECT  3.05 5.55 4.30 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.75 2.50 11.00 ;
        RECT  4.50 7.75 5.20 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 3.65 ;
        RECT  8.65 2.00 10.25 2.70 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.40 4.25 2.10 4.95 ;
        RECT  3.00 3.15 3.50 4.75 ;
        RECT  1.40 4.25 3.50 4.75 ;
        RECT  3.15 6.80 3.85 9.45 ;
        RECT  3.15 6.80 6.55 7.30 ;
        RECT  5.15 2.95 5.85 3.65 ;
        RECT  5.85 6.80 6.55 10.55 ;
        RECT  7.20 6.80 7.90 9.45 ;
        RECT  8.55 7.75 9.25 10.55 ;
        RECT  5.85 10.05 9.25 10.55 ;
        RECT  7.20 6.80 10.60 7.30 ;
        RECT  9.90 6.80 10.60 10.55 ;
        RECT  11.25 6.80 11.95 9.45 ;
        RECT  12.60 7.75 13.30 10.55 ;
        RECT  9.90 10.05 13.30 10.55 ;
        RECT  13.05 2.95 13.75 3.65 ;
        RECT  11.25 6.80 14.70 7.30 ;
        RECT  3.00 3.15 14.70 3.65 ;
        RECT  14.20 3.15 14.70 9.45 ;
        RECT  13.95 6.80 14.70 9.45 ;
    END
END AO333X1
MACRO AO333X2
    CLASS CORE ;
    FOREIGN AO333X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.70 0.95 10.20 ;
        RECT  0.45 2.70 1.15 3.40 ;
        RECT  0.45 7.35 1.15 10.20 ;
        RECT  0.25 9.30 1.15 10.20 ;
        END
    END Q
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  12.85 4.10 13.75 5.00 ;
        END
    END J
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  10.05 4.10 10.95 5.00 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.40 9.55 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 4.10 5.35 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        RECT  3.05 5.55 4.30 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.75 2.50 11.00 ;
        RECT  4.50 7.75 5.20 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 3.65 ;
        RECT  8.65 2.00 10.25 2.70 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.40 4.25 2.10 4.95 ;
        RECT  3.00 3.15 3.50 4.75 ;
        RECT  1.40 4.25 3.50 4.75 ;
        RECT  3.15 6.80 3.85 9.45 ;
        RECT  3.15 6.80 6.55 7.30 ;
        RECT  5.15 2.95 5.85 3.65 ;
        RECT  5.85 6.80 6.55 10.55 ;
        RECT  7.20 6.80 7.90 9.45 ;
        RECT  8.55 7.75 9.25 10.55 ;
        RECT  5.85 10.05 9.25 10.55 ;
        RECT  7.20 6.80 10.60 7.30 ;
        RECT  9.90 6.80 10.60 10.55 ;
        RECT  11.25 6.80 11.95 9.45 ;
        RECT  12.60 7.75 13.30 10.55 ;
        RECT  9.90 10.05 13.30 10.55 ;
        RECT  13.05 2.95 13.75 3.65 ;
        RECT  11.25 6.80 14.70 7.30 ;
        RECT  3.00 3.15 14.70 3.65 ;
        RECT  14.20 3.15 14.70 9.45 ;
        RECT  13.95 6.80 14.70 9.45 ;
    END
END AO333X2
MACRO AO333X4
    CLASS CORE ;
    FOREIGN AO333X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.45 2.30 10.55 ;
        RECT  1.80 2.45 2.50 4.05 ;
        RECT  1.80 7.95 2.55 10.55 ;
        RECT  1.65 9.30 2.55 10.55 ;
        END
    END Q
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  14.25 4.10 15.15 5.00 ;
        END
    END J
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.80 6.30 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  11.45 4.10 12.35 5.00 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.40 9.55 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 4.10 6.75 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        RECT  4.45 5.55 5.80 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 4.20 7.60 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 8.05 1.15 11.00 ;
        RECT  3.15 8.05 3.85 11.00 ;
        RECT  6.00 7.85 6.70 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.85 ;
        RECT  3.15 2.00 3.85 3.85 ;
        RECT  10.15 2.00 11.75 2.70 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.80 4.40 3.50 5.10 ;
        RECT  4.40 3.15 4.90 4.90 ;
        RECT  2.80 4.40 4.90 4.90 ;
        RECT  4.65 6.90 5.35 9.55 ;
        RECT  4.65 6.90 8.05 7.40 ;
        RECT  6.65 2.95 7.35 3.65 ;
        RECT  7.35 6.90 8.05 10.50 ;
        RECT  8.70 6.90 9.40 9.55 ;
        RECT  10.05 7.85 10.75 10.50 ;
        RECT  7.35 10.00 10.75 10.50 ;
        RECT  8.70 6.90 12.10 7.40 ;
        RECT  11.40 6.90 12.10 10.50 ;
        RECT  12.75 6.90 13.45 9.55 ;
        RECT  14.10 7.85 14.80 10.50 ;
        RECT  11.40 10.00 14.80 10.50 ;
        RECT  14.55 2.95 15.25 3.65 ;
        RECT  12.75 6.90 16.15 7.40 ;
        RECT  4.40 3.15 16.15 3.65 ;
        RECT  15.65 3.15 16.15 9.55 ;
        RECT  15.45 6.90 16.15 9.55 ;
    END
END AO333X4
MACRO AO33X1
    CLASS CORE ;
    FOREIGN AO33X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.25 3.40 0.75 10.20 ;
        RECT  0.25 3.40 1.15 4.10 ;
        RECT  0.25 8.05 1.15 10.20 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  10.05 4.10 10.95 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 4.00 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.55 7.60 ;
        RECT  1.65 6.85 2.85 7.60 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.05 2.50 11.00 ;
        RECT  4.50 8.05 5.20 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.95 2.00 2.65 3.90 ;
        RECT  8.65 2.00 9.35 3.90 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.45 4.45 1.95 5.25 ;
        RECT  1.25 4.55 1.95 5.25 ;
        RECT  3.35 7.05 3.85 9.75 ;
        RECT  3.15 8.05 3.85 9.75 ;
        RECT  3.35 7.05 6.55 7.55 ;
        RECT  5.30 3.20 6.00 4.95 ;
        RECT  5.85 7.05 6.55 10.55 ;
        RECT  7.20 7.05 7.90 9.60 ;
        RECT  1.45 4.45 9.10 4.95 ;
        RECT  1.25 4.55 9.10 4.95 ;
        RECT  8.60 4.45 9.10 7.55 ;
        RECT  8.55 8.05 9.25 10.55 ;
        RECT  5.85 10.05 9.25 10.55 ;
        RECT  7.20 7.05 10.60 7.55 ;
        RECT  9.90 7.05 10.60 9.60 ;
    END
END AO33X1
MACRO AO33X2
    CLASS CORE ;
    FOREIGN AO33X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.25 2.50 0.75 10.50 ;
        RECT  0.25 2.50 1.15 4.10 ;
        RECT  0.25 8.00 1.15 10.50 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  10.05 4.10 10.95 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 4.00 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.55 7.60 ;
        RECT  1.65 6.85 2.85 7.60 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.05 2.50 11.00 ;
        RECT  4.50 8.05 5.20 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.00 ;
        RECT  8.65 2.00 9.35 3.90 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.45 4.45 1.95 5.25 ;
        RECT  1.25 4.55 1.95 5.25 ;
        RECT  3.35 7.05 3.85 9.75 ;
        RECT  3.15 8.05 3.85 9.75 ;
        RECT  3.35 7.05 6.55 7.55 ;
        RECT  5.30 3.20 6.00 4.95 ;
        RECT  5.85 7.05 6.55 10.55 ;
        RECT  7.20 7.05 7.90 9.60 ;
        RECT  1.45 4.45 9.10 4.95 ;
        RECT  1.25 4.55 9.10 4.95 ;
        RECT  8.60 4.45 9.10 7.55 ;
        RECT  8.55 8.05 9.25 10.55 ;
        RECT  5.85 10.05 9.25 10.55 ;
        RECT  7.20 7.05 10.60 7.55 ;
        RECT  9.90 7.05 10.60 9.60 ;
    END
END AO33X2
MACRO AO33X4
    CLASS CORE ;
    FOREIGN AO33X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.85 2.50 2.15 10.50 ;
        RECT  1.65 3.60 2.15 10.50 ;
        RECT  1.85 2.50 2.55 4.10 ;
        RECT  1.65 3.60 2.55 4.10 ;
        RECT  1.65 8.00 2.55 10.50 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.40 9.55 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.40 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        RECT  3.05 6.85 4.25 7.60 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 8.05 1.15 11.00 ;
        RECT  3.15 8.05 3.85 11.00 ;
        RECT  6.00 8.05 6.70 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 2.00 1.20 4.00 ;
        RECT  3.20 2.00 3.90 4.00 ;
        RECT  10.05 2.00 10.75 3.90 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.85 4.45 3.35 5.25 ;
        RECT  2.65 4.55 3.35 5.25 ;
        RECT  4.85 7.05 5.35 9.75 ;
        RECT  4.65 8.05 5.35 9.75 ;
        RECT  4.85 7.05 8.05 7.55 ;
        RECT  6.70 3.20 7.40 4.95 ;
        RECT  7.35 7.05 8.05 10.55 ;
        RECT  8.70 7.05 9.40 9.60 ;
        RECT  2.85 4.45 10.50 4.95 ;
        RECT  2.65 4.55 10.50 4.95 ;
        RECT  10.00 4.45 10.50 7.55 ;
        RECT  10.05 8.05 10.75 10.55 ;
        RECT  7.35 10.05 10.75 10.55 ;
        RECT  8.70 7.05 12.10 7.55 ;
        RECT  11.40 7.05 12.10 9.60 ;
    END
END AO33X4
MACRO BTHCX12
    CLASS CORE ;
    FOREIGN BTHCX12 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.65 6.75 9.45 10.55 ;
        RECT  9.60 2.45 10.30 4.60 ;
        RECT  9.80 2.45 10.30 6.30 ;
        RECT  10.40 5.40 10.90 7.25 ;
        RECT  9.80 5.40 10.95 6.30 ;
        RECT  11.35 6.75 12.15 10.55 ;
        RECT  12.75 2.45 13.45 4.60 ;
        RECT  12.95 2.45 13.45 5.90 ;
        RECT  9.80 5.40 13.45 5.90 ;
        RECT  8.65 6.75 14.85 7.25 ;
        RECT  14.05 6.75 14.85 10.55 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.24 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.66 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.95 9.70 3.75 11.00 ;
        RECT  4.60 7.70 5.40 11.00 ;
        RECT  7.30 7.10 8.10 11.00 ;
        RECT  10.00 7.70 10.80 11.00 ;
        RECT  12.70 7.70 13.50 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.20 2.00 2.90 3.25 ;
        RECT  4.90 2.00 5.60 3.25 ;
        RECT  8.25 2.00 8.95 4.50 ;
        RECT  11.40 2.00 11.65 4.45 ;
        RECT  10.95 3.10 11.65 4.45 ;
        RECT  11.40 2.00 12.10 3.55 ;
        RECT  10.95 3.10 12.10 3.55 ;
        RECT  14.25 2.00 14.95 4.50 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.50 2.45 1.30 3.30 ;
        RECT  0.80 2.45 1.30 4.75 ;
        RECT  1.10 6.75 1.60 10.45 ;
        RECT  1.10 8.70 1.80 10.45 ;
        RECT  1.60 4.25 2.10 7.25 ;
        RECT  1.10 6.75 2.10 7.25 ;
        RECT  2.65 4.05 3.35 4.75 ;
        RECT  0.80 4.25 3.35 4.75 ;
        RECT  2.95 6.75 3.75 7.85 ;
        RECT  3.50 2.45 4.30 3.40 ;
        RECT  3.80 2.45 4.30 4.95 ;
        RECT  4.40 4.45 4.90 7.25 ;
        RECT  2.95 6.75 4.90 7.25 ;
        RECT  3.80 4.45 6.30 4.95 ;
        RECT  5.60 4.45 6.30 5.25 ;
        RECT  6.25 5.85 6.75 10.55 ;
        RECT  5.95 7.05 6.75 10.55 ;
        RECT  6.75 3.55 7.50 4.30 ;
        RECT  7.00 3.55 7.50 6.35 ;
        RECT  7.00 5.65 8.40 6.35 ;
        RECT  6.25 5.85 8.40 6.35 ;
    END
END BTHCX12
MACRO BTHCX16
    CLASS CORE ;
    FOREIGN BTHCX16 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.55 6.80 12.35 10.55 ;
        RECT  12.95 2.45 13.65 4.60 ;
        RECT  13.15 2.45 13.65 5.40 ;
        RECT  14.25 6.80 15.05 10.55 ;
        RECT  15.65 2.45 16.40 5.40 ;
        RECT  17.10 6.80 17.90 10.55 ;
        RECT  18.35 2.45 19.10 5.40 ;
        RECT  18.45 2.45 19.10 6.30 ;
        RECT  18.45 5.40 19.35 6.30 ;
        RECT  18.85 2.45 19.10 7.30 ;
        RECT  13.15 4.90 19.10 5.40 ;
        RECT  18.85 5.40 19.35 7.30 ;
        RECT  11.55 6.80 20.60 7.30 ;
        RECT  19.80 6.80 20.60 10.55 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.85 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.32 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.25 7.05 0.75 11.00 ;
        RECT  0.25 10.65 1.60 11.00 ;
        RECT  0.25 7.05 1.65 8.90 ;
        RECT  4.85 7.40 5.60 11.00 ;
        RECT  7.50 7.70 8.30 11.00 ;
        RECT  10.20 7.75 11.00 11.00 ;
        RECT  12.90 7.75 13.70 11.00 ;
        RECT  15.65 7.75 16.50 11.00 ;
        RECT  18.45 7.75 19.25 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.55 2.00 3.25 4.50 ;
        RECT  2.55 2.00 4.45 2.25 ;
        RECT  6.45 2.00 7.15 4.00 ;
        RECT  8.20 2.00 10.75 2.10 ;
        RECT  11.60 2.00 12.30 4.50 ;
        RECT  14.30 2.00 15.00 4.45 ;
        RECT  17.00 2.00 17.70 4.45 ;
        RECT  19.85 2.00 20.55 4.50 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.90 2.95 2.10 3.65 ;
        RECT  1.60 2.95 2.10 5.75 ;
        RECT  1.60 5.05 2.65 5.75 ;
        RECT  2.15 5.05 2.65 10.45 ;
        RECT  2.15 9.65 3.80 10.45 ;
        RECT  3.90 2.80 4.40 8.70 ;
        RECT  3.25 7.10 4.40 8.70 ;
        RECT  3.90 2.80 4.60 4.95 ;
        RECT  5.10 2.55 5.80 3.30 ;
        RECT  3.90 2.80 5.80 3.30 ;
        RECT  6.15 6.75 6.95 10.55 ;
        RECT  3.90 4.45 10.05 4.95 ;
        RECT  8.95 3.30 9.65 4.00 ;
        RECT  9.20 5.85 9.65 10.55 ;
        RECT  8.85 6.75 9.65 10.55 ;
        RECT  9.20 5.85 9.70 7.25 ;
        RECT  6.15 6.75 9.70 7.25 ;
        RECT  9.35 4.45 10.05 5.15 ;
        RECT  8.95 3.50 11.15 4.00 ;
        RECT  10.65 3.50 11.15 6.35 ;
        RECT  10.65 5.65 11.40 6.35 ;
        RECT  9.20 5.85 11.40 6.35 ;
    END
END BTHCX16
MACRO BTHCX20
    CLASS CORE ;
    FOREIGN BTHCX20 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.60 6.80 12.40 10.55 ;
        RECT  12.95 2.45 13.65 4.60 ;
        RECT  13.15 2.45 13.65 5.40 ;
        RECT  14.30 6.80 15.10 10.55 ;
        RECT  15.65 2.45 16.40 5.40 ;
        RECT  17.15 6.80 17.95 10.55 ;
        RECT  18.35 2.45 19.10 5.40 ;
        RECT  18.45 2.45 19.10 6.30 ;
        RECT  18.45 5.40 19.35 6.30 ;
        RECT  18.85 2.45 19.10 7.30 ;
        RECT  13.15 4.90 19.10 5.40 ;
        RECT  18.85 5.40 19.35 7.30 ;
        RECT  11.60 6.80 20.65 7.30 ;
        RECT  19.85 6.80 20.65 10.15 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.85 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.32 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.25 7.10 0.75 11.00 ;
        RECT  0.25 7.10 1.70 8.70 ;
        RECT  0.25 10.70 1.80 11.00 ;
        RECT  4.85 7.40 5.65 11.00 ;
        RECT  7.55 7.70 8.35 11.00 ;
        RECT  10.25 7.20 11.05 11.00 ;
        RECT  12.95 7.75 13.75 11.00 ;
        RECT  15.70 7.75 16.55 11.00 ;
        RECT  18.50 7.75 19.30 11.00 ;
        RECT  21.20 7.10 22.00 11.00 ;
        RECT  0.00 11.00 22.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.55 2.00 3.25 4.50 ;
        RECT  2.55 2.00 4.45 2.25 ;
        RECT  6.45 2.00 7.15 4.00 ;
        RECT  8.20 2.00 10.75 2.10 ;
        RECT  11.60 2.00 12.30 4.50 ;
        RECT  14.30 2.00 15.00 4.45 ;
        RECT  17.00 2.00 17.70 4.45 ;
        RECT  19.70 2.00 20.40 4.45 ;
        RECT  21.25 2.00 21.95 4.50 ;
        RECT  0.00 0.00 22.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.90 2.95 2.10 3.65 ;
        RECT  1.60 2.95 2.10 5.75 ;
        RECT  1.60 5.05 2.70 5.75 ;
        RECT  2.20 5.05 2.70 9.65 ;
        RECT  2.95 9.15 3.55 10.45 ;
        RECT  2.20 9.15 3.55 9.65 ;
        RECT  2.95 9.65 3.65 10.45 ;
        RECT  3.90 2.80 4.40 8.70 ;
        RECT  3.35 7.10 4.40 8.70 ;
        RECT  3.90 2.80 4.60 4.95 ;
        RECT  5.10 2.55 5.80 3.30 ;
        RECT  3.90 2.80 5.80 3.30 ;
        RECT  6.20 6.75 7.00 10.55 ;
        RECT  6.20 6.75 9.70 7.25 ;
        RECT  3.90 4.45 10.05 4.95 ;
        RECT  8.95 3.30 9.65 4.00 ;
        RECT  9.20 5.85 9.70 10.55 ;
        RECT  8.90 6.75 9.70 10.55 ;
        RECT  9.35 4.45 10.05 5.15 ;
        RECT  8.95 3.50 11.15 4.00 ;
        RECT  10.65 3.50 11.15 6.35 ;
        RECT  10.65 5.65 11.45 6.35 ;
        RECT  9.20 5.85 11.45 6.35 ;
    END
END BTHCX20
MACRO BTHCX3
    CLASS CORE ;
    FOREIGN BTHCX3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.90 6.75 9.40 10.55 ;
        RECT  8.60 7.95 9.40 10.55 ;
        RECT  10.00 2.45 10.70 4.60 ;
        RECT  10.25 2.45 10.70 7.25 ;
        RECT  10.20 2.45 10.70 6.30 ;
        RECT  10.25 5.40 10.75 7.25 ;
        RECT  8.90 6.75 10.75 7.25 ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.58 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.48 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.35 7.60 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.40 7.10 1.20 11.00 ;
        RECT  4.40 8.90 5.20 11.00 ;
        RECT  3.30 9.70 5.20 11.00 ;
        RECT  7.25 8.25 8.05 11.00 ;
        RECT  9.95 7.95 10.75 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.30 2.00 2.00 2.60 ;
        RECT  2.75 2.00 3.55 4.25 ;
        RECT  5.45 2.00 6.25 4.40 ;
        RECT  8.65 2.00 9.35 4.50 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.25 3.55 2.30 4.25 ;
        RECT  1.80 3.55 2.30 9.65 ;
        RECT  1.80 7.30 2.50 8.00 ;
        RECT  1.80 4.70 2.65 5.40 ;
        RECT  1.80 8.95 2.85 9.65 ;
        RECT  3.50 5.65 4.00 7.80 ;
        RECT  3.30 7.10 4.00 7.80 ;
        RECT  4.10 3.50 4.90 4.40 ;
        RECT  4.40 3.50 4.90 6.15 ;
        RECT  6.05 7.30 6.55 10.55 ;
        RECT  5.75 8.95 6.55 10.55 ;
        RECT  5.90 5.45 6.60 6.15 ;
        RECT  3.50 5.65 6.60 6.15 ;
        RECT  7.10 3.70 7.90 4.45 ;
        RECT  7.40 3.70 7.90 7.80 ;
        RECT  6.05 7.30 7.90 7.80 ;
        RECT  7.40 6.80 8.45 7.50 ;
        RECT  6.05 7.30 8.45 7.50 ;
    END
END BTHCX3
MACRO BTHCX4
    CLASS CORE ;
    FOREIGN BTHCX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.90 6.75 9.40 10.55 ;
        RECT  8.60 7.95 9.40 10.55 ;
        RECT  9.85 2.45 10.55 4.60 ;
        RECT  10.35 2.45 10.55 7.25 ;
        RECT  10.05 2.45 10.55 6.30 ;
        RECT  10.35 5.40 10.85 7.25 ;
        RECT  8.90 6.75 10.85 7.25 ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.58 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.48 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.35 7.60 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.30 1.15 11.00 ;
        RECT  4.45 8.90 5.15 11.00 ;
        RECT  3.30 9.70 5.15 11.00 ;
        RECT  7.25 7.95 8.05 11.00 ;
        RECT  9.95 7.95 10.75 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.25 2.00 2.00 2.60 ;
        RECT  2.75 2.00 3.55 4.25 ;
        RECT  5.45 2.00 6.25 4.40 ;
        RECT  8.50 2.00 9.20 4.50 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 7.25 2.50 7.95 ;
        RECT  1.25 3.60 2.30 4.40 ;
        RECT  2.00 3.60 2.30 9.65 ;
        RECT  1.80 3.60 2.30 7.95 ;
        RECT  2.00 7.25 2.50 9.65 ;
        RECT  2.00 8.95 2.85 9.65 ;
        RECT  1.80 4.70 3.05 5.40 ;
        RECT  3.50 5.65 4.00 7.80 ;
        RECT  3.30 7.10 4.00 7.80 ;
        RECT  4.10 3.50 4.90 4.40 ;
        RECT  4.40 3.50 4.90 6.15 ;
        RECT  6.05 7.00 6.55 10.55 ;
        RECT  5.75 8.95 6.55 10.55 ;
        RECT  6.05 5.45 6.75 6.15 ;
        RECT  3.50 5.65 6.75 6.15 ;
        RECT  7.00 3.70 7.70 4.45 ;
        RECT  7.20 3.70 7.70 7.50 ;
        RECT  7.20 6.80 8.45 7.50 ;
        RECT  6.05 7.00 8.45 7.50 ;
    END
END BTHCX4
MACRO BTHCX8
    CLASS CORE ;
    FOREIGN BTHCX8 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.65 6.75 9.45 10.55 ;
        RECT  9.60 2.45 10.30 4.60 ;
        RECT  9.80 2.45 10.30 6.30 ;
        RECT  10.40 5.40 10.90 7.25 ;
        RECT  9.80 5.40 10.95 6.30 ;
        RECT  8.65 6.75 12.15 7.25 ;
        RECT  11.35 6.75 12.15 10.55 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.24 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.66 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.95 9.70 3.75 11.00 ;
        RECT  4.60 7.70 5.40 11.00 ;
        RECT  7.30 7.10 8.10 11.00 ;
        RECT  10.00 7.70 10.80 11.00 ;
        RECT  12.70 7.70 13.50 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.20 2.00 2.90 3.25 ;
        RECT  4.90 2.00 5.60 3.25 ;
        RECT  8.25 2.00 8.95 4.50 ;
        RECT  11.30 2.00 12.05 4.45 ;
        RECT  10.95 3.40 12.05 4.45 ;
        RECT  12.85 2.00 13.55 4.50 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.50 2.45 1.30 3.30 ;
        RECT  0.80 2.45 1.30 4.75 ;
        RECT  1.10 6.75 1.60 10.45 ;
        RECT  1.10 8.70 1.80 10.45 ;
        RECT  1.60 4.25 2.10 7.25 ;
        RECT  1.10 6.75 2.10 7.25 ;
        RECT  2.65 4.05 3.35 4.75 ;
        RECT  0.80 4.25 3.35 4.75 ;
        RECT  2.95 6.75 3.75 7.85 ;
        RECT  3.50 2.45 4.30 3.40 ;
        RECT  3.80 2.45 4.30 4.95 ;
        RECT  4.40 4.45 4.90 7.25 ;
        RECT  2.95 6.75 4.90 7.25 ;
        RECT  3.80 4.45 6.30 4.95 ;
        RECT  5.60 4.45 6.30 5.25 ;
        RECT  6.25 5.85 6.75 10.55 ;
        RECT  5.95 7.05 6.75 10.55 ;
        RECT  6.75 3.55 7.50 4.30 ;
        RECT  7.00 3.55 7.50 6.35 ;
        RECT  7.00 5.65 8.40 6.35 ;
        RECT  6.25 5.85 8.40 6.35 ;
    END
END BTHCX8
MACRO BTHX1
    CLASS CORE ;
    FOREIGN BTHX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.50 3.35 9.55 4.05 ;
        RECT  8.65 5.40 9.55 6.30 ;
        RECT  9.05 3.35 9.55 10.10 ;
        RECT  8.65 8.35 9.55 10.10 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.45 1.15 11.00 ;
        RECT  4.45 10.25 5.15 11.00 ;
        RECT  7.30 8.35 8.00 11.00 ;
        RECT  7.15 10.45 8.00 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.75 ;
        RECT  7.15 2.00 7.85 4.00 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.80 5.40 3.80 5.90 ;
        RECT  0.95 3.40 2.10 4.10 ;
        RECT  1.80 3.40 2.10 9.15 ;
        RECT  1.60 3.40 2.10 7.05 ;
        RECT  1.80 6.35 2.50 9.15 ;
        RECT  2.55 3.60 3.30 4.30 ;
        RECT  1.60 6.35 2.85 7.05 ;
        RECT  2.80 3.60 3.30 5.90 ;
        RECT  3.30 5.40 3.80 9.80 ;
        RECT  3.30 7.15 4.00 9.80 ;
        RECT  4.65 2.70 4.80 8.85 ;
        RECT  4.10 2.70 4.80 4.95 ;
        RECT  4.65 4.45 5.15 8.85 ;
        RECT  4.65 7.15 5.35 8.85 ;
        RECT  3.30 9.30 6.50 9.80 ;
        RECT  5.80 3.35 6.50 4.95 ;
        RECT  6.00 7.40 6.50 10.55 ;
        RECT  5.80 9.30 6.50 10.55 ;
        RECT  4.10 4.45 8.25 4.95 ;
        RECT  7.55 4.45 8.25 5.15 ;
        RECT  7.75 7.20 8.45 7.90 ;
        RECT  6.00 7.40 8.45 7.90 ;
    END
END BTHX1
MACRO BTHX12
    CLASS CORE ;
    FOREIGN BTHX12 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.80 2.45 9.50 4.05 ;
        RECT  9.00 2.45 9.50 10.55 ;
        RECT  8.80 7.70 9.50 10.55 ;
        RECT  11.45 2.45 11.95 10.55 ;
        RECT  11.45 2.45 12.20 4.05 ;
        RECT  11.45 7.70 12.20 10.55 ;
        RECT  11.45 5.40 12.35 6.30 ;
        RECT  9.00 5.40 14.70 5.90 ;
        RECT  14.20 2.45 14.70 10.55 ;
        RECT  14.20 2.45 14.90 4.05 ;
        RECT  14.20 7.70 14.90 10.55 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.65 9.25 1.35 11.00 ;
        RECT  4.60 9.95 5.30 11.00 ;
        RECT  7.45 7.70 8.15 11.00 ;
        RECT  10.15 7.25 10.85 11.00 ;
        RECT  12.85 7.25 13.55 11.00 ;
        RECT  15.55 7.25 16.25 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.60 ;
        RECT  7.45 2.00 8.15 4.00 ;
        RECT  10.15 2.00 10.85 4.00 ;
        RECT  12.85 2.00 13.55 4.00 ;
        RECT  15.55 2.00 16.25 4.00 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.60 6.05 2.35 6.75 ;
        RECT  2.80 6.85 3.95 7.35 ;
        RECT  0.95 3.25 2.10 3.95 ;
        RECT  1.85 3.25 2.10 10.45 ;
        RECT  1.60 3.25 2.10 6.75 ;
        RECT  1.85 6.05 2.35 10.45 ;
        RECT  1.85 9.75 2.70 10.45 ;
        RECT  2.55 3.45 3.30 4.15 ;
        RECT  3.25 3.45 3.30 9.50 ;
        RECT  2.80 3.45 3.30 7.35 ;
        RECT  3.25 6.85 3.95 9.50 ;
        RECT  4.10 2.55 4.80 4.95 ;
        RECT  4.80 4.45 5.30 8.55 ;
        RECT  4.60 6.85 5.30 8.55 ;
        RECT  3.25 9.00 6.80 9.50 ;
        RECT  6.10 2.45 6.80 4.95 ;
        RECT  6.30 6.75 6.80 10.55 ;
        RECT  6.10 7.70 6.80 10.55 ;
        RECT  4.10 4.45 8.50 4.95 ;
        RECT  7.80 4.45 8.50 5.15 ;
        RECT  7.85 6.15 8.55 7.25 ;
        RECT  6.30 6.75 8.55 7.25 ;
    END
END BTHX12
MACRO BTHX16
    CLASS CORE ;
    FOREIGN BTHX16 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  9.00 2.45 9.70 4.05 ;
        RECT  9.20 2.45 9.70 10.55 ;
        RECT  9.00 7.70 9.70 10.55 ;
        RECT  11.70 2.45 12.40 4.05 ;
        RECT  11.45 5.40 12.40 6.30 ;
        RECT  11.90 2.45 12.40 10.55 ;
        RECT  11.70 7.70 12.40 10.55 ;
        RECT  14.40 2.45 14.90 10.55 ;
        RECT  14.40 2.45 15.10 4.05 ;
        RECT  14.40 7.70 15.10 10.55 ;
        RECT  9.20 5.40 17.60 5.90 ;
        RECT  17.10 2.45 17.60 10.55 ;
        RECT  17.10 2.45 17.80 4.05 ;
        RECT  17.10 7.70 17.80 10.55 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.65 9.25 1.35 11.00 ;
        RECT  4.55 9.95 5.25 11.00 ;
        RECT  7.65 7.70 8.35 11.00 ;
        RECT  10.35 7.25 11.05 11.00 ;
        RECT  13.05 7.25 13.75 11.00 ;
        RECT  15.75 7.25 16.45 11.00 ;
        RECT  18.45 7.25 19.15 11.00 ;
        RECT  0.00 11.00 19.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.60 ;
        RECT  7.50 2.00 8.20 4.00 ;
        RECT  10.35 2.00 11.05 4.00 ;
        RECT  13.05 2.00 13.75 4.00 ;
        RECT  15.75 2.00 16.45 4.00 ;
        RECT  18.45 2.00 19.15 4.00 ;
        RECT  0.00 0.00 19.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.60 6.05 2.35 6.75 ;
        RECT  2.80 6.85 3.90 7.35 ;
        RECT  0.95 3.25 2.10 3.95 ;
        RECT  1.85 3.25 2.10 10.45 ;
        RECT  1.60 3.25 2.10 6.75 ;
        RECT  1.85 6.05 2.35 10.45 ;
        RECT  1.85 9.75 2.70 10.45 ;
        RECT  2.55 3.45 3.30 4.15 ;
        RECT  3.20 3.45 3.30 9.50 ;
        RECT  2.80 3.45 3.30 7.35 ;
        RECT  3.20 6.85 3.90 9.50 ;
        RECT  4.75 2.55 4.80 8.55 ;
        RECT  4.10 2.55 4.80 4.95 ;
        RECT  4.75 4.45 5.25 8.55 ;
        RECT  4.55 6.85 5.25 8.55 ;
        RECT  3.20 9.00 6.90 9.50 ;
        RECT  6.15 2.45 6.85 4.95 ;
        RECT  6.40 6.75 6.90 10.55 ;
        RECT  6.20 8.05 6.90 10.55 ;
        RECT  4.10 4.45 8.70 4.95 ;
        RECT  8.00 4.45 8.70 5.15 ;
        RECT  8.05 5.70 8.75 7.25 ;
        RECT  6.40 6.75 8.75 7.25 ;
    END
END BTHX16
MACRO BTHX2
    CLASS CORE ;
    FOREIGN BTHX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.65 2.45 9.55 4.05 ;
        RECT  9.05 2.45 9.55 10.55 ;
        RECT  8.65 7.70 9.55 10.55 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.45 1.15 11.00 ;
        RECT  4.45 10.25 5.15 11.00 ;
        RECT  7.30 7.70 8.00 11.00 ;
        RECT  7.15 10.75 8.00 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.75 ;
        RECT  7.30 2.00 8.00 4.00 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.80 5.40 3.80 5.90 ;
        RECT  0.95 3.40 2.10 4.10 ;
        RECT  1.80 3.40 2.10 9.15 ;
        RECT  1.60 3.40 2.10 7.05 ;
        RECT  1.80 6.35 2.50 9.15 ;
        RECT  2.55 3.60 3.30 4.30 ;
        RECT  1.60 6.35 2.85 7.05 ;
        RECT  2.80 3.60 3.30 5.90 ;
        RECT  3.30 5.40 3.80 9.80 ;
        RECT  3.30 7.15 4.00 9.80 ;
        RECT  4.65 2.70 4.80 8.85 ;
        RECT  4.10 2.70 4.80 4.95 ;
        RECT  4.65 4.45 5.15 8.85 ;
        RECT  4.65 7.15 5.35 8.85 ;
        RECT  3.30 9.30 6.50 9.80 ;
        RECT  5.80 3.35 6.50 4.95 ;
        RECT  6.00 6.75 6.50 10.55 ;
        RECT  5.80 9.30 6.50 10.55 ;
        RECT  4.10 4.45 8.40 4.95 ;
        RECT  7.70 4.45 8.40 5.15 ;
        RECT  7.75 6.15 8.45 7.25 ;
        RECT  6.00 6.75 8.45 7.25 ;
    END
END BTHX2
MACRO BTHX20
    CLASS CORE ;
    FOREIGN BTHX20 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  9.10 2.45 9.80 4.05 ;
        RECT  9.30 2.45 9.80 10.55 ;
        RECT  9.10 7.70 9.80 10.55 ;
        RECT  11.80 2.45 12.50 4.05 ;
        RECT  12.00 2.45 12.50 10.55 ;
        RECT  11.80 7.70 12.50 10.55 ;
        RECT  14.50 2.45 15.20 4.05 ;
        RECT  14.25 5.40 15.20 6.30 ;
        RECT  14.70 2.45 15.20 10.55 ;
        RECT  14.50 7.70 15.20 10.55 ;
        RECT  17.20 2.45 17.70 10.55 ;
        RECT  17.20 2.45 17.90 4.05 ;
        RECT  17.20 7.70 17.90 10.55 ;
        RECT  9.30 5.40 20.40 5.90 ;
        RECT  19.90 2.45 20.40 10.55 ;
        RECT  19.90 2.45 20.60 4.05 ;
        RECT  19.90 7.70 20.60 10.55 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.20 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 9.45 1.15 11.00 ;
        RECT  3.35 9.95 4.05 11.00 ;
        RECT  7.75 7.70 8.45 11.00 ;
        RECT  10.45 7.25 11.15 11.00 ;
        RECT  13.15 7.25 13.85 11.00 ;
        RECT  15.85 7.25 16.55 11.00 ;
        RECT  18.55 7.25 19.25 11.00 ;
        RECT  21.25 7.25 21.95 11.00 ;
        RECT  0.00 11.00 22.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.60 ;
        RECT  7.65 2.00 8.35 4.00 ;
        RECT  10.45 2.00 11.15 4.00 ;
        RECT  13.15 2.00 13.85 4.00 ;
        RECT  15.85 2.00 16.55 4.00 ;
        RECT  18.55 2.00 19.25 4.00 ;
        RECT  21.25 2.00 21.95 4.00 ;
        RECT  0.00 0.00 22.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.15 4.45 2.10 4.95 ;
        RECT  0.95 3.25 1.65 3.95 ;
        RECT  1.60 3.25 1.65 10.55 ;
        RECT  1.15 3.25 1.65 4.95 ;
        RECT  1.60 4.45 2.10 10.55 ;
        RECT  1.60 5.60 2.35 6.30 ;
        RECT  1.60 9.85 2.50 10.55 ;
        RECT  2.50 3.45 3.30 4.15 ;
        RECT  2.55 6.85 3.30 8.55 ;
        RECT  2.80 3.45 3.30 9.50 ;
        RECT  4.05 2.55 4.60 8.55 ;
        RECT  3.90 6.85 4.60 8.55 ;
        RECT  2.80 9.00 5.20 9.50 ;
        RECT  4.05 2.55 4.75 4.95 ;
        RECT  4.70 9.00 5.20 10.55 ;
        RECT  5.85 2.45 7.00 3.15 ;
        RECT  5.50 7.90 7.10 8.60 ;
        RECT  6.40 7.90 7.10 10.55 ;
        RECT  6.30 2.45 7.00 4.95 ;
        RECT  6.60 6.75 7.10 10.55 ;
        RECT  4.70 9.85 7.10 10.55 ;
        RECT  4.05 4.45 8.80 4.95 ;
        RECT  8.10 4.45 8.80 5.15 ;
        RECT  8.15 5.70 8.85 7.25 ;
        RECT  6.60 6.75 8.85 7.25 ;
    END
END BTHX20
MACRO BTHX3
    CLASS CORE ;
    FOREIGN BTHX3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.65 3.25 9.55 3.95 ;
        RECT  9.05 3.25 9.55 10.20 ;
        RECT  8.65 7.60 9.55 10.20 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.45 1.15 11.00 ;
        RECT  4.45 10.25 5.15 11.00 ;
        RECT  7.35 7.70 8.05 11.00 ;
        RECT  7.15 9.75 8.05 11.00 ;
        RECT  10.05 7.60 10.75 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.75 ;
        RECT  7.30 2.00 8.00 3.95 ;
        RECT  10.00 2.00 10.70 3.95 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.80 5.40 3.80 5.90 ;
        RECT  0.95 3.40 2.10 4.10 ;
        RECT  1.80 3.40 2.10 9.15 ;
        RECT  1.60 3.40 2.10 7.05 ;
        RECT  1.80 6.35 2.50 9.15 ;
        RECT  2.55 3.60 3.30 4.30 ;
        RECT  1.60 6.35 2.85 7.05 ;
        RECT  2.80 3.60 3.30 5.90 ;
        RECT  3.30 5.40 3.80 9.80 ;
        RECT  3.30 7.15 4.00 9.80 ;
        RECT  4.65 2.70 4.80 8.85 ;
        RECT  4.10 2.70 4.80 4.95 ;
        RECT  4.65 4.45 5.15 8.85 ;
        RECT  4.65 7.15 5.35 8.85 ;
        RECT  3.30 9.30 6.50 9.80 ;
        RECT  5.80 3.50 6.50 4.95 ;
        RECT  6.00 6.75 6.50 10.55 ;
        RECT  5.80 9.30 6.50 10.55 ;
        RECT  4.10 4.45 8.40 4.95 ;
        RECT  7.65 6.25 8.35 7.25 ;
        RECT  6.00 6.75 8.35 7.25 ;
        RECT  7.70 4.45 8.40 5.30 ;
    END
END BTHX3
MACRO BTHX4
    CLASS CORE ;
    FOREIGN BTHX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.65 2.45 9.55 4.05 ;
        RECT  9.05 2.45 9.55 10.55 ;
        RECT  8.70 7.70 9.55 10.55 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.45 1.15 11.00 ;
        RECT  4.45 10.25 5.15 11.00 ;
        RECT  7.30 7.70 8.05 11.00 ;
        RECT  7.15 10.75 8.05 11.00 ;
        RECT  10.05 7.25 10.75 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.75 ;
        RECT  7.35 2.00 8.05 4.00 ;
        RECT  10.05 2.00 10.75 4.00 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.80 5.40 3.80 5.90 ;
        RECT  0.95 3.40 2.10 4.10 ;
        RECT  1.80 3.40 2.10 9.15 ;
        RECT  1.60 3.40 2.10 7.05 ;
        RECT  1.80 6.35 2.50 9.15 ;
        RECT  2.55 3.60 3.30 4.30 ;
        RECT  1.60 6.35 2.85 7.05 ;
        RECT  2.80 3.60 3.30 5.90 ;
        RECT  3.30 5.40 3.80 9.80 ;
        RECT  3.30 7.15 4.00 9.80 ;
        RECT  4.65 2.70 4.80 8.85 ;
        RECT  4.10 2.70 4.80 4.95 ;
        RECT  4.65 4.45 5.15 8.85 ;
        RECT  4.65 7.15 5.35 8.85 ;
        RECT  3.30 9.30 6.50 9.80 ;
        RECT  5.80 3.35 6.50 4.95 ;
        RECT  6.00 6.75 6.50 10.55 ;
        RECT  5.80 9.30 6.50 10.55 ;
        RECT  4.10 4.45 8.40 4.95 ;
        RECT  7.70 4.45 8.40 5.15 ;
        RECT  7.75 6.15 8.45 7.25 ;
        RECT  6.00 6.75 8.45 7.25 ;
    END
END BTHX4
MACRO BTHX8
    CLASS CORE ;
    FOREIGN BTHX8 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.65 2.45 9.55 4.05 ;
        RECT  9.05 2.45 9.55 10.55 ;
        RECT  8.80 7.70 9.55 10.55 ;
        RECT  9.05 5.15 11.90 5.65 ;
        RECT  11.40 2.45 11.90 10.55 ;
        RECT  11.40 2.45 12.10 4.05 ;
        RECT  11.40 7.70 12.20 10.55 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.65 9.25 1.35 11.00 ;
        RECT  4.60 9.95 5.30 11.00 ;
        RECT  7.45 7.70 8.15 11.00 ;
        RECT  10.15 7.25 10.85 11.00 ;
        RECT  12.85 7.25 13.55 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.60 ;
        RECT  7.35 2.00 8.05 4.00 ;
        RECT  10.05 2.00 10.75 4.00 ;
        RECT  12.75 2.00 13.45 4.00 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.60 6.05 2.35 6.75 ;
        RECT  2.80 6.85 3.95 7.35 ;
        RECT  0.95 3.25 2.10 3.95 ;
        RECT  1.85 3.25 2.10 10.45 ;
        RECT  1.60 3.25 2.10 6.75 ;
        RECT  1.85 6.05 2.35 10.45 ;
        RECT  1.85 9.75 2.70 10.45 ;
        RECT  2.55 3.45 3.30 4.15 ;
        RECT  3.25 3.45 3.30 9.50 ;
        RECT  2.80 3.45 3.30 7.35 ;
        RECT  3.25 6.85 3.95 9.50 ;
        RECT  4.10 2.55 4.80 4.95 ;
        RECT  4.80 4.45 5.30 8.55 ;
        RECT  4.60 6.85 5.30 8.55 ;
        RECT  3.25 9.00 6.80 9.50 ;
        RECT  6.00 2.45 6.70 4.95 ;
        RECT  6.10 6.75 6.80 10.55 ;
        RECT  4.10 4.45 8.40 4.95 ;
        RECT  7.70 4.45 8.40 5.15 ;
        RECT  7.90 6.15 8.60 7.25 ;
        RECT  6.10 6.75 8.60 7.25 ;
    END
END BTHX8
MACRO BTLCX12
    CLASS CORE ;
    FOREIGN BTLCX12 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.05 6.75 10.85 10.55 ;
        RECT  10.90 2.45 11.60 4.60 ;
        RECT  11.45 2.45 11.60 7.25 ;
        RECT  11.10 2.45 11.60 5.90 ;
        RECT  11.45 5.40 12.30 7.25 ;
        RECT  11.45 5.40 12.35 6.30 ;
        RECT  12.75 6.75 13.55 10.55 ;
        RECT  13.60 3.55 14.30 4.50 ;
        RECT  13.80 3.55 14.30 5.90 ;
        RECT  14.10 2.45 14.30 5.90 ;
        RECT  11.10 5.40 14.30 5.90 ;
        RECT  14.10 2.45 14.80 4.05 ;
        RECT  13.60 3.55 14.80 4.05 ;
        RECT  15.45 6.75 16.25 10.55 ;
        RECT  10.05 6.75 16.30 7.25 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.68 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.35 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.66 ;
        PORT
        LAYER M1M ;
        RECT  2.95 5.40 3.95 6.45 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 7.90 1.25 11.00 ;
        RECT  4.55 9.20 5.25 11.00 ;
        RECT  6.05 7.70 6.80 11.00 ;
        RECT  8.70 7.10 9.50 11.00 ;
        RECT  11.40 7.70 12.20 11.00 ;
        RECT  14.10 7.70 14.90 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.45 2.00 4.30 4.45 ;
        RECT  6.30 2.00 7.00 3.25 ;
        RECT  9.55 2.00 10.25 4.50 ;
        RECT  12.70 2.00 13.00 4.45 ;
        RECT  12.25 2.60 13.00 4.45 ;
        RECT  12.70 2.00 13.45 3.00 ;
        RECT  12.25 2.60 13.45 3.00 ;
        RECT  15.65 2.00 16.35 4.50 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.75 2.50 2.50 4.55 ;
        RECT  2.00 2.50 2.50 8.40 ;
        RECT  2.00 7.30 2.60 8.40 ;
        RECT  1.90 7.70 2.60 8.40 ;
        RECT  2.00 7.30 4.45 7.80 ;
        RECT  3.25 8.25 3.75 10.35 ;
        RECT  3.05 9.15 3.75 10.35 ;
        RECT  3.75 7.10 4.45 7.80 ;
        RECT  1.90 7.70 4.45 7.80 ;
        RECT  4.90 2.55 5.40 8.75 ;
        RECT  3.25 8.25 5.40 8.75 ;
        RECT  4.90 2.55 5.65 3.25 ;
        RECT  4.90 4.45 7.60 4.95 ;
        RECT  6.90 4.45 7.60 5.20 ;
        RECT  7.65 5.85 8.15 10.55 ;
        RECT  7.35 7.05 8.15 10.55 ;
        RECT  8.05 3.55 8.90 4.25 ;
        RECT  8.40 3.55 8.90 6.35 ;
        RECT  8.40 5.65 9.80 6.35 ;
        RECT  7.65 5.85 9.80 6.35 ;
    END
END BTLCX12
MACRO BTLCX16
    CLASS CORE ;
    FOREIGN BTLCX16 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.55 6.80 12.35 10.55 ;
        RECT  12.95 2.45 13.65 4.60 ;
        RECT  13.15 2.45 13.65 5.40 ;
        RECT  14.25 6.80 15.05 10.55 ;
        RECT  15.65 2.45 16.40 5.40 ;
        RECT  17.10 6.80 17.90 10.55 ;
        RECT  18.35 2.45 19.10 5.40 ;
        RECT  18.45 2.45 19.10 7.30 ;
        RECT  13.15 4.90 19.10 5.40 ;
        RECT  18.45 5.40 19.35 7.30 ;
        RECT  11.55 6.80 20.60 7.30 ;
        RECT  19.80 6.80 20.60 10.55 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.73 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.35 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.32 ;
        PORT
        LAYER M1M ;
        RECT  5.80 5.40 6.75 6.35 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.90 7.20 1.70 11.00 ;
        RECT  4.85 7.40 5.60 11.00 ;
        RECT  7.50 7.75 8.30 11.00 ;
        RECT  10.20 7.75 11.00 11.00 ;
        RECT  12.90 7.75 13.70 11.00 ;
        RECT  15.65 7.75 16.50 11.00 ;
        RECT  18.45 7.75 19.25 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.55 2.00 3.25 4.40 ;
        RECT  2.55 2.00 4.45 2.25 ;
        RECT  6.45 2.00 7.15 4.00 ;
        RECT  8.20 2.00 10.75 2.10 ;
        RECT  11.60 2.00 12.30 4.50 ;
        RECT  14.30 2.00 15.00 4.45 ;
        RECT  17.00 2.00 17.70 4.45 ;
        RECT  19.85 2.00 20.55 4.50 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.70 2.50 1.40 3.20 ;
        RECT  0.90 2.50 1.40 4.25 ;
        RECT  0.90 3.55 2.10 4.25 ;
        RECT  1.60 3.55 2.10 5.35 ;
        RECT  1.60 4.85 2.65 5.35 ;
        RECT  2.15 4.85 2.65 10.55 ;
        RECT  2.15 9.85 4.30 10.55 ;
        RECT  3.90 2.80 4.40 8.85 ;
        RECT  3.25 7.25 4.40 8.85 ;
        RECT  3.90 2.80 4.60 4.95 ;
        RECT  5.10 2.55 5.80 3.30 ;
        RECT  3.90 2.80 5.80 3.30 ;
        RECT  6.15 6.80 6.95 10.55 ;
        RECT  3.90 4.45 10.05 4.95 ;
        RECT  8.95 3.30 9.65 4.00 ;
        RECT  9.20 5.85 9.65 10.55 ;
        RECT  8.85 6.80 9.65 10.55 ;
        RECT  9.20 5.85 9.70 7.30 ;
        RECT  6.15 6.80 9.70 7.30 ;
        RECT  9.35 4.45 10.05 5.15 ;
        RECT  8.95 3.50 11.15 4.00 ;
        RECT  10.65 3.50 11.15 6.35 ;
        RECT  10.65 5.65 11.40 6.35 ;
        RECT  9.20 5.85 11.40 6.35 ;
    END
END BTLCX16
MACRO BTLCX20
    CLASS CORE ;
    FOREIGN BTLCX20 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.55 6.80 12.35 10.55 ;
        RECT  12.95 2.45 13.65 4.60 ;
        RECT  13.15 2.45 13.65 5.40 ;
        RECT  14.25 6.80 15.05 10.55 ;
        RECT  15.65 2.45 16.40 5.40 ;
        RECT  16.95 6.80 17.75 10.55 ;
        RECT  18.35 2.45 19.10 5.40 ;
        RECT  18.45 2.45 19.10 6.30 ;
        RECT  18.45 5.40 19.35 6.30 ;
        RECT  18.85 2.45 19.10 7.30 ;
        RECT  13.15 4.90 19.10 5.40 ;
        RECT  18.85 5.40 19.35 7.30 ;
        RECT  11.55 6.80 20.45 7.30 ;
        RECT  19.65 6.80 20.45 10.55 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.73 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.32 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 7.20 1.65 11.00 ;
        RECT  4.85 7.40 5.60 11.00 ;
        RECT  7.50 7.70 8.30 11.00 ;
        RECT  10.20 7.75 11.00 11.00 ;
        RECT  12.90 7.75 13.70 11.00 ;
        RECT  15.65 7.75 16.35 11.00 ;
        RECT  18.30 7.75 19.10 11.00 ;
        RECT  21.15 6.90 21.95 11.00 ;
        RECT  0.00 11.00 22.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.55 2.00 3.25 4.40 ;
        RECT  2.55 2.00 4.45 2.25 ;
        RECT  6.45 2.00 7.15 4.00 ;
        RECT  8.20 2.00 10.75 2.10 ;
        RECT  11.60 2.00 12.30 4.50 ;
        RECT  14.30 2.00 15.00 4.45 ;
        RECT  17.00 2.00 17.70 4.45 ;
        RECT  19.70 2.00 20.40 4.55 ;
        RECT  21.25 2.00 21.95 4.50 ;
        RECT  0.00 0.00 22.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.70 2.45 1.40 3.15 ;
        RECT  0.90 2.45 1.40 4.25 ;
        RECT  0.90 3.55 2.10 4.25 ;
        RECT  1.60 3.55 2.10 5.45 ;
        RECT  1.60 4.85 2.65 5.45 ;
        RECT  2.15 4.85 2.65 10.55 ;
        RECT  2.15 9.80 4.35 10.55 ;
        RECT  3.90 2.80 4.40 8.85 ;
        RECT  3.25 7.25 4.40 8.85 ;
        RECT  3.90 2.80 4.60 4.95 ;
        RECT  5.10 2.55 5.80 3.30 ;
        RECT  3.90 2.80 5.80 3.30 ;
        RECT  6.15 6.75 6.95 10.55 ;
        RECT  3.90 4.45 10.05 4.95 ;
        RECT  8.95 3.30 9.65 4.00 ;
        RECT  9.20 5.85 9.65 10.55 ;
        RECT  8.85 6.75 9.65 10.55 ;
        RECT  9.20 5.85 9.70 7.25 ;
        RECT  6.15 6.75 9.70 7.25 ;
        RECT  9.35 4.45 10.05 5.15 ;
        RECT  8.95 3.50 11.15 4.00 ;
        RECT  10.65 3.50 11.15 6.35 ;
        RECT  10.65 5.65 11.40 6.35 ;
        RECT  9.20 5.85 11.40 6.35 ;
    END
END BTLCX20
MACRO BTLCX3
    CLASS CORE ;
    FOREIGN BTLCX3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.90 6.75 9.40 10.55 ;
        RECT  8.60 7.95 9.40 10.55 ;
        RECT  10.00 2.45 10.70 4.60 ;
        RECT  10.25 2.45 10.70 7.25 ;
        RECT  10.20 2.45 10.70 6.30 ;
        RECT  10.25 5.40 10.75 7.25 ;
        RECT  8.90 6.75 10.75 7.25 ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.16 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.48 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.40 7.10 1.20 11.00 ;
        RECT  0.40 10.05 2.50 11.00 ;
        RECT  4.40 9.20 5.20 11.00 ;
        RECT  3.30 9.70 5.20 11.00 ;
        RECT  7.30 8.25 8.05 11.00 ;
        RECT  9.95 7.95 10.75 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 2.00 3.55 4.25 ;
        RECT  5.45 2.00 6.25 4.25 ;
        RECT  8.65 2.00 9.35 4.50 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.95 2.60 1.65 3.30 ;
        RECT  1.15 2.60 1.65 4.35 ;
        RECT  1.15 3.65 2.30 4.35 ;
        RECT  1.80 3.65 2.30 8.75 ;
        RECT  1.80 7.30 2.50 8.75 ;
        RECT  3.30 6.80 4.00 7.80 ;
        RECT  4.10 3.50 4.90 4.70 ;
        RECT  4.40 3.50 4.90 7.30 ;
        RECT  3.30 6.80 4.90 7.30 ;
        RECT  4.70 7.80 5.20 8.75 ;
        RECT  1.80 8.25 5.20 8.75 ;
        RECT  4.40 4.70 6.60 5.20 ;
        RECT  4.70 7.80 5.90 8.50 ;
        RECT  1.80 8.25 5.90 8.50 ;
        RECT  5.90 4.70 6.60 5.40 ;
        RECT  6.35 7.30 6.85 10.55 ;
        RECT  5.75 8.95 6.85 10.55 ;
        RECT  7.10 3.70 7.90 4.45 ;
        RECT  7.40 3.70 7.90 7.80 ;
        RECT  6.35 7.30 7.90 7.80 ;
        RECT  7.40 6.80 8.45 7.50 ;
        RECT  6.35 7.30 8.45 7.50 ;
    END
END BTLCX3
MACRO BTLCX4
    CLASS CORE ;
    FOREIGN BTLCX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.90 5.80 9.40 10.55 ;
        RECT  8.65 7.10 9.40 10.55 ;
        RECT  9.85 2.45 10.55 4.60 ;
        RECT  10.05 2.45 10.55 6.30 ;
        RECT  10.05 5.40 10.95 6.30 ;
        RECT  8.90 5.80 10.95 6.30 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.16 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.48 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.40 7.10 1.20 11.00 ;
        RECT  0.40 10.05 2.50 11.00 ;
        RECT  4.45 9.20 5.15 11.00 ;
        RECT  3.35 9.75 5.15 11.00 ;
        RECT  7.30 7.10 8.00 11.00 ;
        RECT  10.00 7.10 10.70 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 2.00 3.55 4.25 ;
        RECT  5.45 2.00 6.25 4.25 ;
        RECT  8.50 2.00 9.20 4.50 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.95 2.60 1.65 3.30 ;
        RECT  1.15 2.60 1.65 4.35 ;
        RECT  1.15 3.65 2.30 4.35 ;
        RECT  1.80 3.65 2.30 8.75 ;
        RECT  1.80 7.30 2.50 8.75 ;
        RECT  3.30 6.80 4.00 7.80 ;
        RECT  4.10 3.50 4.90 4.70 ;
        RECT  4.40 3.50 4.90 7.30 ;
        RECT  3.30 6.80 4.90 7.30 ;
        RECT  4.70 7.80 5.20 8.75 ;
        RECT  1.80 8.25 5.20 8.75 ;
        RECT  4.40 4.70 6.60 5.20 ;
        RECT  4.70 7.80 5.90 8.50 ;
        RECT  1.80 8.25 5.90 8.50 ;
        RECT  6.35 6.15 6.50 10.55 ;
        RECT  5.80 8.95 6.50 10.55 ;
        RECT  5.90 4.70 6.60 5.40 ;
        RECT  6.35 6.15 6.85 9.45 ;
        RECT  5.80 8.95 6.85 9.45 ;
        RECT  6.95 3.70 7.90 4.40 ;
        RECT  7.40 3.70 7.90 6.65 ;
        RECT  7.40 5.95 8.45 6.65 ;
        RECT  6.35 6.15 8.45 6.65 ;
    END
END BTLCX4
MACRO BTLCX8
    CLASS CORE ;
    FOREIGN BTLCX8 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.05 6.75 10.85 10.55 ;
        RECT  11.00 2.45 11.70 4.60 ;
        RECT  11.50 2.45 11.70 7.25 ;
        RECT  11.20 2.45 11.70 6.30 ;
        RECT  11.50 5.40 12.30 7.25 ;
        RECT  11.20 5.40 12.35 6.30 ;
        RECT  10.05 6.75 13.55 7.25 ;
        RECT  12.75 6.75 13.55 10.55 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.68 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.35 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.66 ;
        PORT
        LAYER M1M ;
        RECT  2.95 5.40 3.95 6.45 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 7.90 1.25 11.00 ;
        RECT  4.55 9.20 5.25 11.00 ;
        RECT  6.05 7.70 6.80 11.00 ;
        RECT  8.70 7.10 9.50 11.00 ;
        RECT  11.40 7.70 12.20 11.00 ;
        RECT  14.10 7.15 14.90 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.45 2.00 4.30 4.45 ;
        RECT  6.30 2.00 7.00 3.25 ;
        RECT  9.65 2.00 10.35 4.50 ;
        RECT  12.70 2.00 13.45 4.45 ;
        RECT  12.35 3.40 13.45 4.45 ;
        RECT  14.25 2.00 14.95 4.50 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.75 2.50 2.50 4.55 ;
        RECT  2.00 2.50 2.50 8.40 ;
        RECT  2.00 7.30 2.60 8.40 ;
        RECT  1.90 7.70 2.60 8.40 ;
        RECT  2.00 7.30 4.45 7.80 ;
        RECT  3.25 8.25 3.75 10.35 ;
        RECT  3.05 9.65 3.75 10.35 ;
        RECT  3.75 7.10 4.45 7.80 ;
        RECT  1.90 7.70 4.45 7.80 ;
        RECT  4.90 2.55 5.40 8.75 ;
        RECT  3.25 8.25 5.40 8.75 ;
        RECT  4.90 2.55 5.65 3.25 ;
        RECT  4.90 4.45 7.70 4.95 ;
        RECT  7.00 4.45 7.70 5.20 ;
        RECT  7.65 5.85 8.15 10.55 ;
        RECT  7.35 7.05 8.15 10.55 ;
        RECT  8.15 3.55 8.90 4.25 ;
        RECT  8.40 3.55 8.90 6.35 ;
        RECT  8.40 5.65 9.80 6.35 ;
        RECT  7.65 5.85 9.80 6.35 ;
    END
END BTLCX8
MACRO BTLX1
    CLASS CORE ;
    FOREIGN BTLX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.50 2.80 9.55 4.05 ;
        RECT  9.05 2.80 9.55 10.10 ;
        RECT  8.65 8.35 9.55 10.10 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.45 1.15 11.00 ;
        RECT  4.45 10.25 5.15 11.00 ;
        RECT  7.30 8.35 8.00 11.00 ;
        RECT  7.15 10.75 8.00 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.75 ;
        RECT  7.15 2.00 7.85 4.00 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.60 4.70 2.30 5.40 ;
        RECT  2.80 5.40 3.80 5.90 ;
        RECT  1.80 3.40 2.10 9.15 ;
        RECT  1.80 7.45 2.50 9.15 ;
        RECT  0.95 3.40 2.10 4.10 ;
        RECT  2.00 3.40 2.10 10.55 ;
        RECT  1.60 3.40 2.10 5.40 ;
        RECT  2.00 4.70 2.30 10.55 ;
        RECT  1.80 4.70 2.30 9.15 ;
        RECT  2.00 7.45 2.50 10.55 ;
        RECT  2.55 3.60 3.30 4.30 ;
        RECT  2.00 9.85 2.85 10.55 ;
        RECT  2.80 3.60 3.30 5.90 ;
        RECT  3.30 5.40 3.80 9.80 ;
        RECT  3.30 7.15 4.00 9.80 ;
        RECT  4.65 2.70 4.80 8.85 ;
        RECT  4.10 2.70 4.80 4.95 ;
        RECT  4.65 4.45 5.15 8.85 ;
        RECT  4.65 7.15 5.35 8.85 ;
        RECT  3.30 9.30 6.50 9.80 ;
        RECT  5.80 3.35 6.50 4.95 ;
        RECT  6.00 7.40 6.50 10.55 ;
        RECT  5.80 9.30 6.50 10.55 ;
        RECT  4.10 4.45 8.25 4.95 ;
        RECT  7.55 4.45 8.25 5.15 ;
        RECT  7.75 7.20 8.45 7.90 ;
        RECT  6.00 7.40 8.45 7.90 ;
    END
END BTLX1
MACRO BTLX12
    CLASS CORE ;
    FOREIGN BTLX12 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.80 2.45 9.50 4.05 ;
        RECT  9.00 2.45 9.50 10.55 ;
        RECT  8.80 7.70 9.50 10.55 ;
        RECT  11.45 2.45 11.95 10.55 ;
        RECT  11.45 2.45 12.20 4.05 ;
        RECT  11.45 7.70 12.20 10.55 ;
        RECT  11.45 5.40 12.35 6.30 ;
        RECT  9.00 5.40 14.70 5.90 ;
        RECT  14.20 2.45 14.70 10.55 ;
        RECT  14.20 2.45 14.90 4.05 ;
        RECT  14.20 7.70 14.90 10.55 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.65 9.25 1.35 11.00 ;
        RECT  4.60 9.95 5.30 11.00 ;
        RECT  7.45 7.70 8.15 11.00 ;
        RECT  10.15 7.25 10.85 11.00 ;
        RECT  12.85 7.25 13.55 11.00 ;
        RECT  15.55 7.25 16.25 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.60 ;
        RECT  7.45 2.00 8.15 4.00 ;
        RECT  10.15 2.00 10.85 4.00 ;
        RECT  12.85 2.00 13.55 4.00 ;
        RECT  15.55 2.00 16.25 4.00 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.80 6.85 3.95 7.35 ;
        RECT  1.60 7.85 2.50 8.35 ;
        RECT  0.95 3.25 2.10 3.95 ;
        RECT  1.40 3.25 2.10 5.00 ;
        RECT  2.00 3.25 2.10 10.45 ;
        RECT  1.60 3.25 2.10 8.35 ;
        RECT  2.00 7.85 2.50 10.45 ;
        RECT  2.00 9.75 2.70 10.45 ;
        RECT  2.55 3.45 3.30 4.15 ;
        RECT  3.25 3.45 3.30 9.40 ;
        RECT  2.80 3.45 3.30 7.35 ;
        RECT  2.00 9.85 4.15 10.45 ;
        RECT  3.25 6.85 3.95 9.40 ;
        RECT  3.45 9.85 4.15 10.55 ;
        RECT  4.10 2.55 4.80 4.95 ;
        RECT  4.80 4.45 5.30 8.45 ;
        RECT  4.60 6.85 5.30 8.45 ;
        RECT  3.25 8.90 6.80 9.40 ;
        RECT  6.10 2.45 6.80 4.95 ;
        RECT  6.30 6.75 6.80 10.55 ;
        RECT  6.10 7.70 6.80 10.55 ;
        RECT  4.10 4.45 8.50 4.95 ;
        RECT  7.80 4.45 8.50 5.15 ;
        RECT  7.85 6.15 8.55 7.25 ;
        RECT  6.30 6.75 8.55 7.25 ;
    END
END BTLX12
MACRO BTLX16
    CLASS CORE ;
    FOREIGN BTLX16 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  9.00 2.45 9.70 4.05 ;
        RECT  9.20 2.45 9.70 10.55 ;
        RECT  9.00 7.70 9.70 10.55 ;
        RECT  11.70 2.45 12.40 4.05 ;
        RECT  11.45 5.40 12.40 6.30 ;
        RECT  11.90 2.45 12.40 10.55 ;
        RECT  11.70 7.70 12.40 10.55 ;
        RECT  14.40 2.45 14.90 10.55 ;
        RECT  14.40 2.45 15.10 4.05 ;
        RECT  14.40 7.70 15.10 10.55 ;
        RECT  9.20 5.40 17.60 5.90 ;
        RECT  17.10 2.45 17.60 10.55 ;
        RECT  17.10 2.45 17.80 4.05 ;
        RECT  17.10 7.70 17.80 10.55 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.65 9.25 1.35 11.00 ;
        RECT  4.55 9.95 5.25 11.00 ;
        RECT  7.65 7.70 8.35 11.00 ;
        RECT  10.35 7.25 11.05 11.00 ;
        RECT  13.05 7.25 13.75 11.00 ;
        RECT  15.75 7.25 16.45 11.00 ;
        RECT  18.45 7.25 19.15 11.00 ;
        RECT  0.00 11.00 19.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.60 ;
        RECT  7.50 2.00 8.20 4.00 ;
        RECT  10.35 2.00 11.05 4.00 ;
        RECT  13.05 2.00 13.75 4.00 ;
        RECT  15.75 2.00 16.45 4.00 ;
        RECT  18.45 2.00 19.15 4.00 ;
        RECT  0.00 0.00 19.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.80 6.85 3.90 7.35 ;
        RECT  1.60 7.80 2.50 8.30 ;
        RECT  0.95 3.25 2.10 3.95 ;
        RECT  1.40 3.25 2.10 5.00 ;
        RECT  2.00 3.25 2.10 10.45 ;
        RECT  1.60 3.25 2.10 8.30 ;
        RECT  2.00 7.80 2.50 10.45 ;
        RECT  2.00 9.75 2.70 10.45 ;
        RECT  2.55 3.45 3.30 4.15 ;
        RECT  3.20 3.45 3.30 9.40 ;
        RECT  2.80 3.45 3.30 7.35 ;
        RECT  2.00 9.85 4.10 10.45 ;
        RECT  3.20 6.85 3.90 9.40 ;
        RECT  3.40 9.85 4.10 10.55 ;
        RECT  4.75 2.55 4.80 8.45 ;
        RECT  4.10 2.55 4.80 4.95 ;
        RECT  4.75 4.45 5.25 8.45 ;
        RECT  4.55 6.85 5.25 8.45 ;
        RECT  3.20 8.90 6.90 9.40 ;
        RECT  6.15 2.45 6.85 4.95 ;
        RECT  6.40 6.75 6.90 10.55 ;
        RECT  6.20 8.05 6.90 10.55 ;
        RECT  4.10 4.45 8.70 4.95 ;
        RECT  8.00 4.45 8.70 5.15 ;
        RECT  8.05 5.70 8.75 7.25 ;
        RECT  6.40 6.75 8.75 7.25 ;
    END
END BTLX16
MACRO BTLX2
    CLASS CORE ;
    FOREIGN BTLX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.65 2.45 9.55 4.05 ;
        RECT  9.05 2.45 9.55 10.55 ;
        RECT  8.65 7.70 9.55 10.55 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.45 1.15 11.00 ;
        RECT  4.45 10.25 5.15 11.00 ;
        RECT  7.30 7.70 8.00 11.00 ;
        RECT  7.15 10.75 8.00 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.75 ;
        RECT  7.30 2.00 8.00 4.00 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.60 4.70 2.30 5.40 ;
        RECT  2.80 5.40 3.80 5.90 ;
        RECT  1.80 3.40 2.10 9.15 ;
        RECT  1.80 7.45 2.50 9.15 ;
        RECT  0.95 3.40 2.10 4.10 ;
        RECT  2.00 3.40 2.10 10.55 ;
        RECT  1.60 3.40 2.10 5.40 ;
        RECT  2.00 4.70 2.30 10.55 ;
        RECT  1.80 4.70 2.30 9.15 ;
        RECT  2.00 7.45 2.50 10.55 ;
        RECT  2.55 3.60 3.30 4.30 ;
        RECT  2.00 9.85 2.85 10.55 ;
        RECT  2.80 3.60 3.30 5.90 ;
        RECT  3.30 5.40 3.80 9.80 ;
        RECT  3.30 7.15 4.00 9.80 ;
        RECT  4.65 2.70 4.80 8.85 ;
        RECT  4.10 2.70 4.80 4.95 ;
        RECT  4.65 4.45 5.15 8.85 ;
        RECT  4.65 7.15 5.35 8.85 ;
        RECT  3.30 9.30 6.50 9.80 ;
        RECT  5.80 3.35 6.50 4.95 ;
        RECT  6.00 6.75 6.50 10.55 ;
        RECT  5.80 9.30 6.50 10.55 ;
        RECT  4.10 4.45 8.40 4.95 ;
        RECT  7.70 4.45 8.40 5.15 ;
        RECT  7.75 6.15 8.45 7.25 ;
        RECT  6.00 6.75 8.45 7.25 ;
    END
END BTLX2
MACRO BTLX20
    CLASS CORE ;
    FOREIGN BTLX20 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  9.10 2.45 9.80 4.05 ;
        RECT  9.30 2.45 9.80 10.55 ;
        RECT  9.10 7.70 9.80 10.55 ;
        RECT  11.80 2.45 12.50 4.05 ;
        RECT  12.00 2.45 12.50 10.55 ;
        RECT  11.80 7.70 12.50 10.55 ;
        RECT  14.50 2.45 15.20 4.05 ;
        RECT  14.25 5.40 15.20 6.30 ;
        RECT  14.70 2.45 15.20 10.55 ;
        RECT  14.50 7.70 15.20 10.55 ;
        RECT  17.20 2.45 17.70 10.55 ;
        RECT  17.20 2.45 17.90 4.05 ;
        RECT  17.20 7.70 17.90 10.55 ;
        RECT  9.30 5.40 20.40 5.90 ;
        RECT  19.90 2.45 20.40 10.55 ;
        RECT  19.90 2.45 20.60 4.05 ;
        RECT  19.90 7.70 20.60 10.55 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.20 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 9.90 1.15 11.00 ;
        RECT  3.35 9.95 4.05 11.00 ;
        RECT  7.75 7.70 8.45 11.00 ;
        RECT  10.45 7.25 11.15 11.00 ;
        RECT  13.15 7.25 13.85 11.00 ;
        RECT  15.85 7.25 16.55 11.00 ;
        RECT  18.55 7.25 19.25 11.00 ;
        RECT  21.25 7.25 21.95 11.00 ;
        RECT  0.00 11.00 22.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.50 ;
        RECT  7.65 2.00 8.35 4.00 ;
        RECT  10.45 2.00 11.15 4.00 ;
        RECT  13.15 2.00 13.85 4.00 ;
        RECT  15.85 2.00 16.55 4.00 ;
        RECT  18.55 2.00 19.25 4.00 ;
        RECT  21.25 2.00 21.95 4.00 ;
        RECT  0.00 0.00 22.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.40 4.20 2.10 4.90 ;
        RECT  0.95 3.15 1.90 3.85 ;
        RECT  1.40 7.95 2.10 8.65 ;
        RECT  1.60 3.15 1.90 10.55 ;
        RECT  1.40 3.15 1.90 4.90 ;
        RECT  1.60 4.20 2.10 10.55 ;
        RECT  1.60 9.85 2.50 10.55 ;
        RECT  2.50 2.95 3.25 3.65 ;
        RECT  2.55 6.45 3.25 8.05 ;
        RECT  2.75 2.95 3.25 9.45 ;
        RECT  4.05 2.45 4.60 8.25 ;
        RECT  3.90 6.65 4.60 8.25 ;
        RECT  2.75 8.95 5.20 9.45 ;
        RECT  4.05 2.45 4.75 3.15 ;
        RECT  4.70 8.95 5.20 10.55 ;
        RECT  5.85 2.45 7.00 3.15 ;
        RECT  5.50 7.90 7.10 8.60 ;
        RECT  6.40 7.90 7.10 10.55 ;
        RECT  6.30 2.45 7.00 4.95 ;
        RECT  6.60 6.75 7.10 10.55 ;
        RECT  4.70 9.85 7.10 10.55 ;
        RECT  4.05 4.45 8.80 4.95 ;
        RECT  8.10 4.45 8.80 5.15 ;
        RECT  8.15 5.70 8.85 7.25 ;
        RECT  6.60 6.75 8.85 7.25 ;
    END
END BTLX20
MACRO BTLX3
    CLASS CORE ;
    FOREIGN BTLX3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.65 3.20 9.55 3.95 ;
        RECT  9.05 3.20 9.55 10.20 ;
        RECT  8.65 7.60 9.55 10.20 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.45 1.15 11.00 ;
        RECT  4.45 10.25 5.15 11.00 ;
        RECT  7.35 7.70 8.05 11.00 ;
        RECT  7.15 9.70 8.05 11.00 ;
        RECT  10.05 7.60 10.75 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.75 ;
        RECT  7.30 2.00 8.00 3.95 ;
        RECT  10.00 2.00 10.70 3.95 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.60 4.70 2.30 5.40 ;
        RECT  2.80 5.40 3.80 5.90 ;
        RECT  1.80 3.40 2.10 9.15 ;
        RECT  1.80 7.45 2.50 9.15 ;
        RECT  0.95 3.40 2.10 4.10 ;
        RECT  2.00 3.40 2.10 10.55 ;
        RECT  1.60 3.40 2.10 5.40 ;
        RECT  2.00 4.70 2.30 10.55 ;
        RECT  1.80 4.70 2.30 9.15 ;
        RECT  2.00 7.45 2.50 10.55 ;
        RECT  2.55 3.60 3.30 4.30 ;
        RECT  2.00 9.85 2.85 10.55 ;
        RECT  2.80 3.60 3.30 5.90 ;
        RECT  3.30 5.40 3.80 9.80 ;
        RECT  3.30 7.15 4.00 9.80 ;
        RECT  4.65 2.70 4.80 8.85 ;
        RECT  4.10 2.70 4.80 4.95 ;
        RECT  4.65 4.45 5.15 8.85 ;
        RECT  4.65 7.15 5.35 8.85 ;
        RECT  3.30 9.30 6.50 9.80 ;
        RECT  5.80 3.50 6.50 4.95 ;
        RECT  6.00 6.75 6.50 10.55 ;
        RECT  5.80 9.30 6.50 10.55 ;
        RECT  4.10 4.45 8.40 4.95 ;
        RECT  7.65 6.25 8.35 7.25 ;
        RECT  6.00 6.75 8.35 7.25 ;
        RECT  7.70 4.45 8.40 5.30 ;
    END
END BTLX3
MACRO BTLX4
    CLASS CORE ;
    FOREIGN BTLX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.65 2.45 9.55 4.05 ;
        RECT  9.05 2.45 9.55 10.55 ;
        RECT  8.70 7.70 9.55 10.55 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.45 1.15 11.00 ;
        RECT  4.45 10.25 5.15 11.00 ;
        RECT  7.35 7.70 8.05 11.00 ;
        RECT  7.15 10.75 8.05 11.00 ;
        RECT  10.05 7.20 10.75 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.75 ;
        RECT  7.35 2.00 8.05 4.00 ;
        RECT  10.05 2.00 10.75 4.00 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.60 4.70 2.30 5.40 ;
        RECT  2.80 5.40 3.80 5.90 ;
        RECT  1.80 3.40 2.10 9.15 ;
        RECT  1.80 7.45 2.50 9.15 ;
        RECT  0.95 3.40 2.10 4.10 ;
        RECT  2.00 3.40 2.10 10.55 ;
        RECT  1.60 3.40 2.10 5.40 ;
        RECT  2.00 4.70 2.30 10.55 ;
        RECT  1.80 4.70 2.30 9.15 ;
        RECT  2.00 7.45 2.50 10.55 ;
        RECT  2.55 3.60 3.30 4.30 ;
        RECT  2.00 9.85 2.85 10.55 ;
        RECT  2.80 3.60 3.30 5.90 ;
        RECT  3.30 5.40 3.80 9.80 ;
        RECT  3.30 7.15 4.00 9.80 ;
        RECT  4.65 2.70 4.80 8.85 ;
        RECT  4.10 2.70 4.80 4.95 ;
        RECT  4.65 4.45 5.15 8.85 ;
        RECT  4.65 7.15 5.35 8.85 ;
        RECT  3.30 9.30 6.50 9.80 ;
        RECT  5.80 3.35 6.50 4.95 ;
        RECT  6.00 6.75 6.50 10.55 ;
        RECT  5.80 9.30 6.50 10.55 ;
        RECT  4.10 4.45 8.40 4.95 ;
        RECT  7.70 4.45 8.40 5.15 ;
        RECT  7.75 6.15 8.45 7.25 ;
        RECT  6.00 6.75 8.45 7.25 ;
    END
END BTLX4
MACRO BTLX8
    CLASS CORE ;
    FOREIGN BTLX8 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.65 2.45 9.55 4.05 ;
        RECT  9.05 2.45 9.55 10.55 ;
        RECT  8.80 7.70 9.55 10.55 ;
        RECT  9.05 5.15 11.90 5.65 ;
        RECT  11.40 2.45 11.90 10.55 ;
        RECT  11.40 2.45 12.10 4.05 ;
        RECT  11.40 7.70 12.20 10.55 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.65 9.25 1.35 11.00 ;
        RECT  4.60 9.95 5.30 11.00 ;
        RECT  7.45 7.70 8.15 11.00 ;
        RECT  10.15 7.25 10.85 11.00 ;
        RECT  12.85 7.25 13.55 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.60 ;
        RECT  7.35 2.00 8.05 4.00 ;
        RECT  10.05 2.00 10.75 4.00 ;
        RECT  12.75 2.00 13.45 4.00 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.80 6.85 3.95 7.35 ;
        RECT  1.60 7.80 2.50 8.30 ;
        RECT  0.95 3.25 2.10 3.95 ;
        RECT  1.40 3.25 2.10 5.00 ;
        RECT  2.00 3.25 2.10 10.45 ;
        RECT  1.60 3.25 2.10 8.30 ;
        RECT  2.00 7.80 2.50 10.45 ;
        RECT  2.00 9.75 2.70 10.45 ;
        RECT  2.55 3.45 3.30 4.15 ;
        RECT  3.25 3.45 3.30 9.40 ;
        RECT  2.80 3.45 3.30 7.35 ;
        RECT  2.00 9.85 4.15 10.45 ;
        RECT  3.25 6.85 3.95 9.40 ;
        RECT  3.45 9.85 4.15 10.55 ;
        RECT  4.10 2.55 4.80 4.95 ;
        RECT  4.80 4.45 5.30 8.45 ;
        RECT  4.60 6.85 5.30 8.45 ;
        RECT  3.25 8.90 6.80 9.40 ;
        RECT  6.00 2.45 6.70 4.95 ;
        RECT  6.30 6.75 6.80 10.55 ;
        RECT  6.10 7.70 6.80 10.55 ;
        RECT  4.10 4.45 8.40 4.95 ;
        RECT  7.70 4.45 8.40 5.15 ;
        RECT  7.90 6.15 8.60 7.25 ;
        RECT  6.30 6.75 8.60 7.25 ;
    END
END BTLX8
MACRO BUCX12
    CLASS CORE ;
    FOREIGN BUCX12 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  6.75 4.40 10.75 4.60 ;
        RECT  4.60 7.00 5.40 10.55 ;
        RECT  4.60 7.00 8.10 7.50 ;
        RECT  6.95 2.45 7.45 4.90 ;
        RECT  6.75 2.45 7.45 4.60 ;
        RECT  7.60 5.80 8.10 10.55 ;
        RECT  7.30 7.00 8.10 10.55 ;
        RECT  10.05 2.45 10.75 4.90 ;
        RECT  6.95 4.40 10.75 4.90 ;
        RECT  10.25 2.45 10.50 10.55 ;
        RECT  10.00 5.80 10.50 10.55 ;
        RECT  10.25 2.45 10.75 6.30 ;
        RECT  10.00 7.10 10.80 10.55 ;
        RECT  10.05 5.40 10.95 6.30 ;
        RECT  7.60 5.80 10.95 6.30 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.01 ;
        PORT
        LAYER M1M ;
        RECT  0.25 2.80 1.15 3.70 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.55 9.10 1.35 11.00 ;
        RECT  3.25 7.00 4.05 11.00 ;
        RECT  5.95 7.95 6.75 11.00 ;
        RECT  8.65 7.10 9.45 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.40 2.00 3.10 2.70 ;
        RECT  5.40 2.00 6.10 4.30 ;
        RECT  8.70 2.00 8.80 3.95 ;
        RECT  8.10 2.95 8.80 3.95 ;
        RECT  8.70 2.00 9.40 3.45 ;
        RECT  8.10 2.95 9.40 3.45 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.25 4.95 0.75 8.65 ;
        RECT  0.25 8.15 2.70 8.65 ;
        RECT  1.40 4.85 2.10 5.60 ;
        RECT  1.90 6.05 2.40 7.70 ;
        RECT  1.60 6.95 2.40 7.70 ;
        RECT  2.40 3.65 3.10 4.35 ;
        RECT  1.90 8.15 2.70 10.55 ;
        RECT  2.60 3.65 3.10 5.45 ;
        RECT  0.25 4.95 3.10 5.45 ;
        RECT  4.00 2.45 4.75 4.30 ;
        RECT  4.25 2.45 4.75 6.55 ;
        RECT  1.90 6.05 4.75 6.55 ;
        RECT  4.25 5.25 6.55 5.75 ;
        RECT  5.85 5.15 6.55 5.85 ;
    END
END BUCX12
MACRO BUCX16
    CLASS CORE ;
    FOREIGN BUCX16 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  6.10 7.00 6.90 10.55 ;
        RECT  7.70 2.45 8.40 4.70 ;
        RECT  6.10 7.00 9.60 7.50 ;
        RECT  9.10 5.50 9.60 10.55 ;
        RECT  8.80 7.00 9.60 10.55 ;
        RECT  10.40 2.45 11.10 4.70 ;
        RECT  7.70 4.20 11.10 4.70 ;
        RECT  10.60 2.45 11.10 6.00 ;
        RECT  11.40 5.40 12.00 10.55 ;
        RECT  11.40 7.10 12.30 10.55 ;
        RECT  11.40 5.40 12.35 6.30 ;
        RECT  13.10 2.45 13.60 6.00 ;
        RECT  10.60 5.40 13.60 6.00 ;
        RECT  13.10 2.45 13.80 4.70 ;
        RECT  10.60 5.45 14.70 6.00 ;
        RECT  9.10 5.50 14.70 6.00 ;
        RECT  14.20 5.45 14.70 10.55 ;
        RECT  14.20 7.10 15.00 10.55 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.83 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.90 9.25 2.70 11.00 ;
        RECT  4.75 7.10 5.55 11.00 ;
        RECT  7.45 7.95 8.25 11.00 ;
        RECT  10.15 7.10 10.95 11.00 ;
        RECT  12.85 7.10 13.65 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.40 2.00 1.20 4.40 ;
        RECT  0.40 2.00 2.70 2.75 ;
        RECT  3.45 2.00 4.25 4.45 ;
        RECT  6.35 2.00 7.05 4.45 ;
        RECT  9.05 2.00 9.75 3.75 ;
        RECT  11.75 2.00 12.45 4.45 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.55 8.30 1.35 10.55 ;
        RECT  1.95 3.65 2.65 4.40 ;
        RECT  2.15 3.65 2.65 8.80 ;
        RECT  2.15 5.60 3.00 6.30 ;
        RECT  0.55 8.30 4.05 8.80 ;
        RECT  3.45 5.25 3.95 7.80 ;
        RECT  3.15 7.05 3.95 7.80 ;
        RECT  3.25 8.30 4.05 10.55 ;
        RECT  4.80 2.55 5.55 4.45 ;
        RECT  5.05 2.55 5.55 5.75 ;
        RECT  3.45 5.25 7.50 5.75 ;
        RECT  6.80 5.20 7.50 5.90 ;
    END
END BUCX16
MACRO BUCX20
    CLASS CORE ;
    FOREIGN BUCX20 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  6.10 7.00 6.90 10.55 ;
        RECT  7.70 2.45 8.40 4.70 ;
        RECT  6.10 7.00 9.60 7.50 ;
        RECT  9.10 5.45 9.60 10.55 ;
        RECT  8.80 7.00 9.60 10.55 ;
        RECT  10.40 2.45 11.10 4.70 ;
        RECT  7.70 4.20 11.10 4.70 ;
        RECT  10.60 2.45 11.10 5.95 ;
        RECT  11.40 5.40 12.00 10.55 ;
        RECT  11.40 7.10 12.30 10.55 ;
        RECT  11.40 5.40 12.35 6.30 ;
        RECT  13.10 2.45 13.60 5.95 ;
        RECT  10.60 5.40 13.60 5.95 ;
        RECT  13.10 2.45 13.80 4.70 ;
        RECT  9.10 5.45 15.00 5.95 ;
        RECT  14.50 5.45 15.00 10.55 ;
        RECT  14.20 7.10 15.00 10.55 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.83 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.90 9.25 2.70 11.00 ;
        RECT  4.75 7.10 5.55 11.00 ;
        RECT  7.45 7.95 8.25 11.00 ;
        RECT  10.15 7.10 10.95 11.00 ;
        RECT  12.85 7.10 13.65 11.00 ;
        RECT  15.55 7.10 16.35 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.40 2.00 1.25 4.40 ;
        RECT  0.40 2.00 2.75 2.75 ;
        RECT  3.45 2.00 4.25 4.45 ;
        RECT  6.35 2.00 7.05 4.35 ;
        RECT  9.05 2.00 9.75 3.75 ;
        RECT  11.75 2.00 12.45 4.45 ;
        RECT  14.45 2.00 15.15 4.45 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.55 8.30 1.35 10.55 ;
        RECT  2.15 3.65 2.65 8.80 ;
        RECT  2.00 3.65 2.70 4.40 ;
        RECT  2.15 5.60 3.00 6.30 ;
        RECT  0.55 8.30 4.05 8.80 ;
        RECT  3.45 5.25 3.95 7.80 ;
        RECT  3.15 7.05 3.95 7.80 ;
        RECT  3.25 8.30 4.05 10.55 ;
        RECT  4.80 2.55 5.55 4.45 ;
        RECT  5.05 2.55 5.55 5.75 ;
        RECT  3.45 5.25 7.50 5.75 ;
        RECT  6.80 5.20 7.50 5.90 ;
    END
END BUCX20
MACRO BUCX3
    CLASS CORE ;
    FOREIGN BUCX3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.45 7.10 6.55 7.95 ;
        RECT  5.85 2.45 6.55 4.60 ;
        RECT  6.05 2.45 6.55 10.55 ;
        RECT  5.75 7.10 6.55 10.55 ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.95 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.40 7.05 1.20 11.00 ;
        RECT  0.40 7.05 1.35 8.95 ;
        RECT  4.40 8.50 5.20 11.00 ;
        RECT  0.00 11.00 7.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.75 2.45 ;
        RECT  2.60 2.00 3.60 2.45 ;
        RECT  4.50 2.00 5.20 4.50 ;
        RECT  0.00 0.00 7.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.95 4.55 2.50 4.95 ;
        RECT  1.70 3.75 2.15 5.70 ;
        RECT  1.70 4.55 2.50 5.70 ;
        RECT  1.90 3.75 2.15 8.95 ;
        RECT  0.95 3.75 2.15 4.95 ;
        RECT  1.90 4.55 2.50 8.95 ;
        RECT  1.90 7.05 2.70 8.95 ;
        RECT  3.15 3.75 3.65 10.45 ;
        RECT  2.70 9.65 3.65 10.45 ;
        RECT  2.95 3.75 3.75 4.55 ;
        RECT  3.15 5.35 5.40 5.85 ;
        RECT  4.70 5.30 5.40 6.00 ;
    END
END BUCX3
MACRO BUCX4
    CLASS CORE ;
    FOREIGN BUCX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  5.85 2.70 6.55 4.60 ;
        RECT  5.85 5.40 6.35 10.55 ;
        RECT  6.05 2.70 6.35 10.55 ;
        RECT  5.55 7.10 6.35 10.55 ;
        RECT  6.05 2.70 6.55 6.30 ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.95 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.40 7.05 1.20 11.00 ;
        RECT  0.40 7.05 1.35 8.95 ;
        RECT  4.20 7.10 5.00 11.00 ;
        RECT  6.90 7.10 7.70 11.00 ;
        RECT  0.00 11.00 8.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.90 2.00 1.70 2.35 ;
        RECT  2.55 2.00 3.70 2.65 ;
        RECT  4.50 2.00 5.20 4.50 ;
        RECT  7.20 2.00 7.90 4.50 ;
        RECT  0.00 0.00 8.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.90 4.05 2.20 4.55 ;
        RECT  1.70 4.95 2.60 5.75 ;
        RECT  0.90 3.70 1.70 4.55 ;
        RECT  1.90 4.05 2.20 8.95 ;
        RECT  1.70 4.05 2.20 5.75 ;
        RECT  1.90 4.95 2.60 8.95 ;
        RECT  1.90 7.05 2.70 8.95 ;
        RECT  3.15 3.65 3.65 10.45 ;
        RECT  2.70 9.65 3.65 10.45 ;
        RECT  2.90 3.65 3.80 4.50 ;
        RECT  3.15 5.35 5.40 5.85 ;
        RECT  4.70 5.25 5.40 5.95 ;
    END
END BUCX4
MACRO BUCX8
    CLASS CORE ;
    FOREIGN BUCX8 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  5.70 2.70 6.40 4.60 ;
        RECT  5.90 2.70 6.10 10.55 ;
        RECT  5.30 9.60 6.10 10.55 ;
        RECT  5.90 2.70 6.40 10.10 ;
        RECT  5.90 7.10 6.70 10.10 ;
        RECT  5.30 9.60 6.70 10.10 ;
        RECT  5.85 5.40 6.75 6.30 ;
        RECT  7.00 2.45 7.80 3.20 ;
        RECT  5.70 2.70 7.80 3.20 ;
        RECT  5.85 5.80 9.10 6.30 ;
        RECT  8.60 5.80 9.10 10.55 ;
        RECT  8.60 7.10 9.40 10.55 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.01 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.70 7.70 2.55 9.15 ;
        RECT  1.70 8.65 4.75 9.15 ;
        RECT  3.95 8.65 4.75 11.00 ;
        RECT  7.25 7.10 8.05 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.85 2.00 1.65 2.75 ;
        RECT  4.35 2.00 5.05 4.50 ;
        RECT  4.35 2.00 6.45 2.20 ;
        RECT  8.40 2.00 9.10 4.50 ;
        RECT  6.95 3.70 9.10 4.50 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.40 6.75 1.20 10.55 ;
        RECT  0.85 3.65 1.65 4.45 ;
        RECT  0.85 3.95 2.20 4.45 ;
        RECT  1.70 3.95 2.20 7.25 ;
        RECT  1.70 5.65 2.60 7.25 ;
        RECT  0.40 6.75 2.60 7.25 ;
        RECT  2.75 2.45 3.65 4.50 ;
        RECT  0.40 9.75 3.40 10.55 ;
        RECT  3.30 2.45 3.65 7.90 ;
        RECT  3.15 2.45 3.65 5.85 ;
        RECT  3.30 5.35 3.80 7.90 ;
        RECT  3.30 7.10 4.20 7.90 ;
        RECT  3.15 5.35 5.40 5.85 ;
        RECT  4.70 5.25 5.40 5.95 ;
    END
END BUCX8
MACRO BUX1
    CLASS CORE ;
    FOREIGN BUX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  3.15 3.75 3.85 4.45 ;
        RECT  3.35 3.75 3.85 9.70 ;
        RECT  3.05 8.00 3.95 9.70 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.45 5.40 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.05 2.50 11.00 ;
        RECT  0.00 11.00 5.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.45 ;
        RECT  0.00 0.00 5.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.75 0.95 9.70 ;
        RECT  0.45 3.75 1.15 4.45 ;
        RECT  0.45 7.00 1.15 9.70 ;
        RECT  2.20 6.80 2.90 7.50 ;
        RECT  0.45 7.00 2.90 7.50 ;
    END
END BUX1
MACRO BUX12
    CLASS CORE ;
    FOREIGN BUX12 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  3.20 2.45 3.90 4.05 ;
        RECT  3.40 2.45 3.90 10.55 ;
        RECT  3.20 7.45 3.90 10.55 ;
        RECT  5.85 2.45 6.35 10.55 ;
        RECT  5.85 2.45 6.60 4.05 ;
        RECT  5.85 7.45 6.60 10.55 ;
        RECT  5.85 5.30 6.75 6.30 ;
        RECT  3.40 5.30 9.10 5.80 ;
        RECT  8.60 2.45 9.10 10.55 ;
        RECT  8.60 2.45 9.30 4.05 ;
        RECT  8.60 7.45 9.30 10.55 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 7.70 2.55 11.00 ;
        RECT  4.55 7.30 5.25 11.00 ;
        RECT  7.25 7.30 7.95 11.00 ;
        RECT  9.95 7.30 10.65 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 2.00 2.55 4.00 ;
        RECT  4.55 2.00 5.25 4.00 ;
        RECT  7.25 2.00 7.95 4.00 ;
        RECT  9.95 2.00 10.65 4.00 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.50 2.45 1.20 4.95 ;
        RECT  0.50 6.75 1.20 10.55 ;
        RECT  0.50 4.45 2.10 4.95 ;
        RECT  1.60 4.45 2.10 7.25 ;
        RECT  0.50 6.75 2.10 7.25 ;
        RECT  1.60 5.50 2.95 6.20 ;
    END
END BUX12
MACRO BUX16
    CLASS CORE ;
    FOREIGN BUX16 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.70 2.45 5.40 4.05 ;
        RECT  4.90 2.45 5.40 10.55 ;
        RECT  4.70 7.45 5.40 10.55 ;
        RECT  7.40 2.45 8.15 4.05 ;
        RECT  7.25 5.30 8.15 6.30 ;
        RECT  7.65 2.45 8.15 10.55 ;
        RECT  7.40 7.45 8.15 10.55 ;
        RECT  10.10 2.45 10.60 10.55 ;
        RECT  10.10 2.45 10.80 4.05 ;
        RECT  10.10 7.45 10.80 10.55 ;
        RECT  4.90 5.30 13.30 5.80 ;
        RECT  12.80 2.45 13.30 10.55 ;
        RECT  12.80 2.45 13.50 4.05 ;
        RECT  12.80 7.45 13.50 10.55 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 7.30 1.20 11.00 ;
        RECT  3.35 7.70 4.05 11.00 ;
        RECT  6.05 7.30 6.75 11.00 ;
        RECT  8.75 7.30 9.45 11.00 ;
        RECT  11.45 7.30 12.15 11.00 ;
        RECT  14.15 7.30 14.85 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 2.00 1.20 3.90 ;
        RECT  3.35 2.00 4.05 4.00 ;
        RECT  6.05 2.00 6.75 4.00 ;
        RECT  8.75 2.00 9.45 4.00 ;
        RECT  11.45 2.00 12.15 4.00 ;
        RECT  14.15 2.00 14.85 4.00 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.85 3.20 2.55 4.95 ;
        RECT  1.85 6.75 2.55 9.95 ;
        RECT  1.85 4.45 3.60 4.95 ;
        RECT  3.10 4.45 3.60 7.25 ;
        RECT  1.85 6.75 3.60 7.25 ;
        RECT  3.10 5.50 4.45 6.20 ;
    END
END BUX16
MACRO BUX2
    CLASS CORE ;
    FOREIGN BUX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  3.30 2.45 4.00 4.05 ;
        RECT  3.50 2.45 4.00 10.20 ;
        RECT  3.30 7.30 4.00 10.20 ;
        RECT  3.30 2.80 5.35 3.70 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 10.10 1.15 11.00 ;
        RECT  1.95 7.70 2.65 11.00 ;
        RECT  0.00 11.00 5.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.95 2.00 2.65 4.00 ;
        RECT  0.00 0.00 5.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.30 1.15 4.95 ;
        RECT  0.45 6.75 1.15 8.95 ;
        RECT  0.45 4.45 2.10 4.95 ;
        RECT  1.60 4.45 2.10 7.25 ;
        RECT  0.45 6.75 2.10 7.25 ;
        RECT  1.60 5.50 3.05 6.20 ;
    END
END BUX2
MACRO BUX20
    CLASS CORE ;
    FOREIGN BUX20 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.70 2.45 5.40 4.05 ;
        RECT  4.90 2.45 5.40 10.55 ;
        RECT  4.70 7.45 5.40 10.55 ;
        RECT  7.40 2.45 8.15 4.05 ;
        RECT  7.65 2.45 8.15 10.55 ;
        RECT  7.40 7.45 8.15 10.55 ;
        RECT  10.10 2.45 10.60 10.55 ;
        RECT  10.10 2.45 10.80 4.05 ;
        RECT  10.10 7.45 10.80 10.55 ;
        RECT  10.05 5.30 10.95 6.30 ;
        RECT  12.80 2.45 13.30 10.55 ;
        RECT  12.80 2.45 13.50 4.05 ;
        RECT  12.80 7.45 13.50 10.55 ;
        RECT  4.90 5.30 16.00 5.80 ;
        RECT  15.50 2.45 16.00 10.55 ;
        RECT  15.50 2.45 16.20 4.05 ;
        RECT  15.50 7.45 16.20 10.55 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.20 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.65 7.30 1.35 11.00 ;
        RECT  3.35 7.70 4.05 11.00 ;
        RECT  6.05 7.30 6.75 11.00 ;
        RECT  8.75 7.30 9.45 11.00 ;
        RECT  11.45 7.30 12.15 11.00 ;
        RECT  14.15 7.30 14.85 11.00 ;
        RECT  16.85 7.30 17.55 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.65 2.00 1.35 4.00 ;
        RECT  3.35 2.00 4.05 4.00 ;
        RECT  6.05 2.00 6.75 4.00 ;
        RECT  8.75 2.00 9.45 4.00 ;
        RECT  11.45 2.00 12.15 4.00 ;
        RECT  14.15 2.00 14.85 4.00 ;
        RECT  16.85 2.00 17.55 4.00 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.00 2.45 2.70 4.95 ;
        RECT  2.00 6.75 2.70 10.55 ;
        RECT  2.00 4.45 3.60 4.95 ;
        RECT  3.10 4.45 3.60 7.25 ;
        RECT  2.00 6.75 3.60 7.25 ;
        RECT  3.10 5.50 4.45 6.20 ;
    END
END BUX20
MACRO BUX3
    CLASS CORE ;
    FOREIGN BUX3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.70 2.80 5.20 10.05 ;
        RECT  4.50 7.45 5.20 10.05 ;
        RECT  4.45 2.80 5.35 4.20 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 10.10 2.05 11.00 ;
        RECT  3.15 7.50 3.85 11.00 ;
        RECT  5.85 7.50 6.55 11.00 ;
        RECT  0.00 11.00 7.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 2.90 ;
        RECT  3.15 2.00 3.85 4.00 ;
        RECT  5.85 2.00 6.55 4.00 ;
        RECT  0.00 0.00 7.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.70 4.85 4.25 4.95 ;
        RECT  0.70 4.45 1.20 7.90 ;
        RECT  0.70 7.40 2.35 7.90 ;
        RECT  1.65 3.75 2.35 4.95 ;
        RECT  1.65 7.40 2.35 9.05 ;
        RECT  3.55 4.45 4.05 5.55 ;
        RECT  0.70 4.45 4.05 4.95 ;
        RECT  3.55 4.85 4.25 5.55 ;
    END
END BUX3
MACRO BUX4
    CLASS CORE ;
    FOREIGN BUX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.70 2.45 5.20 10.55 ;
        RECT  4.50 7.45 5.20 10.55 ;
        RECT  4.45 2.45 5.35 4.05 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 10.10 2.05 11.00 ;
        RECT  3.15 7.30 3.85 11.00 ;
        RECT  5.85 7.30 6.55 11.00 ;
        RECT  0.00 11.00 7.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.15 2.00 3.85 4.00 ;
        RECT  5.85 2.00 6.55 4.00 ;
        RECT  0.00 0.00 7.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.70 4.55 4.25 4.95 ;
        RECT  0.70 4.45 1.20 7.80 ;
        RECT  0.70 7.30 2.35 7.80 ;
        RECT  1.65 3.50 2.35 4.95 ;
        RECT  1.65 7.30 2.35 8.95 ;
        RECT  3.55 4.45 4.05 5.25 ;
        RECT  0.70 4.45 4.05 4.95 ;
        RECT  3.55 4.55 4.25 5.25 ;
    END
END BUX4
MACRO BUX8
    CLASS CORE ;
    FOREIGN BUX8 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  3.20 2.45 3.90 4.05 ;
        RECT  3.40 2.45 3.90 10.55 ;
        RECT  3.20 7.45 3.90 10.55 ;
        RECT  3.40 5.30 6.75 5.80 ;
        RECT  5.85 2.45 6.35 10.55 ;
        RECT  5.85 2.45 6.60 4.05 ;
        RECT  5.85 7.45 6.60 10.55 ;
        RECT  5.85 5.30 6.75 6.30 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 7.70 2.55 11.00 ;
        RECT  4.55 7.30 5.25 11.00 ;
        RECT  7.25 7.30 7.95 11.00 ;
        RECT  0.00 11.00 8.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 2.00 2.55 4.00 ;
        RECT  4.55 2.00 5.25 4.00 ;
        RECT  7.25 2.00 7.95 4.00 ;
        RECT  0.00 0.00 8.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.50 2.45 1.20 4.95 ;
        RECT  0.50 6.75 1.20 10.55 ;
        RECT  0.50 4.45 2.10 4.95 ;
        RECT  1.60 4.45 2.10 7.25 ;
        RECT  0.50 6.75 2.10 7.25 ;
        RECT  1.60 5.50 2.95 6.20 ;
    END
END BUX8
MACRO DFFRSX1
    CLASS CORE ;
    FOREIGN DFFRSX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 28.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  13.45 5.75 14.15 6.45 ;
        RECT  15.65 5.35 16.55 6.35 ;
        RECT  13.45 5.85 16.55 6.35 ;
        RECT  15.65 5.50 17.75 6.20 ;
        RECT  13.45 5.85 17.75 6.20 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  9.50 2.70 10.95 3.45 ;
        RECT  10.50 2.60 10.95 3.70 ;
        RECT  10.05 2.70 10.95 3.70 ;
        RECT  10.50 2.60 22.50 3.10 ;
        RECT  9.50 2.70 22.50 3.10 ;
        RECT  21.80 2.60 22.50 3.30 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  26.85 2.65 27.35 9.75 ;
        RECT  26.85 2.65 27.55 3.40 ;
        RECT  26.85 8.10 27.55 9.75 ;
        RECT  26.85 5.40 27.75 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  24.15 2.65 24.85 4.30 ;
        RECT  24.15 7.25 24.85 9.75 ;
        RECT  24.15 3.80 25.95 4.30 ;
        RECT  25.45 3.80 25.95 7.75 ;
        RECT  24.15 7.25 25.95 7.75 ;
        RECT  25.45 5.40 26.35 6.30 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.35 7.60 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.40 2.50 11.00 ;
        RECT  4.05 8.05 4.75 11.00 ;
        RECT  3.60 10.75 6.10 11.00 ;
        RECT  9.80 8.30 10.50 11.00 ;
        RECT  12.65 7.30 13.35 11.00 ;
        RECT  12.65 7.30 18.20 7.80 ;
        RECT  17.50 7.30 18.20 8.35 ;
        RECT  19.85 9.25 20.55 11.00 ;
        RECT  22.55 9.25 23.25 11.00 ;
        RECT  25.50 8.25 26.20 11.00 ;
        RECT  0.00 11.00 28.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.20 ;
        RECT  4.05 2.00 4.75 4.85 ;
        RECT  8.50 2.00 9.00 4.95 ;
        RECT  9.90 4.45 10.60 5.20 ;
        RECT  11.45 3.55 11.95 4.95 ;
        RECT  8.50 4.45 11.95 4.95 ;
        RECT  11.45 3.55 14.85 4.05 ;
        RECT  14.15 3.55 14.85 4.25 ;
        RECT  19.85 3.55 20.55 4.25 ;
        RECT  19.85 3.75 23.65 4.25 ;
        RECT  23.15 2.00 23.65 5.50 ;
        RECT  23.15 4.80 24.40 5.50 ;
        RECT  25.50 2.00 26.20 3.30 ;
        RECT  0.00 0.00 28.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.65 3.70 1.15 10.15 ;
        RECT  0.45 9.45 1.15 10.15 ;
        RECT  1.65 5.55 2.60 6.25 ;
        RECT  1.75 2.45 2.25 4.20 ;
        RECT  0.65 3.70 2.25 4.20 ;
        RECT  2.10 5.55 2.60 8.75 ;
        RECT  2.70 4.20 3.40 6.05 ;
        RECT  2.10 8.05 3.40 8.75 ;
        RECT  1.75 2.45 3.55 3.15 ;
        RECT  1.65 5.55 6.35 6.05 ;
        RECT  5.35 3.20 5.85 6.05 ;
        RECT  5.85 5.55 6.35 7.45 ;
        RECT  5.85 6.75 6.55 7.45 ;
        RECT  6.40 4.20 7.55 4.90 ;
        RECT  7.05 4.20 7.55 9.00 ;
        RECT  7.05 3.00 7.75 3.70 ;
        RECT  5.35 3.20 7.75 3.70 ;
        RECT  6.40 8.30 8.15 9.00 ;
        RECT  9.35 5.65 10.05 6.35 ;
        RECT  10.35 6.90 11.05 7.60 ;
        RECT  7.05 7.10 11.05 7.60 ;
        RECT  11.65 5.65 12.15 9.00 ;
        RECT  11.15 8.30 12.15 9.00 ;
        RECT  12.45 4.55 12.95 6.15 ;
        RECT  9.35 5.65 12.95 6.15 ;
        RECT  12.45 4.55 13.15 5.25 ;
        RECT  15.00 8.30 15.70 10.05 ;
        RECT  16.50 3.55 17.20 4.25 ;
        RECT  17.50 8.85 18.20 9.95 ;
        RECT  16.50 3.75 19.35 4.25 ;
        RECT  18.85 3.75 19.35 9.35 ;
        RECT  15.00 8.85 19.35 9.35 ;
        RECT  19.85 4.75 22.05 5.45 ;
        RECT  21.20 8.25 21.90 9.90 ;
        RECT  21.55 4.75 22.05 6.55 ;
        RECT  21.95 7.05 22.65 7.75 ;
        RECT  18.85 7.25 22.65 7.75 ;
        RECT  23.15 6.05 23.65 8.75 ;
        RECT  21.20 8.25 23.65 8.75 ;
        RECT  21.55 6.05 24.95 6.55 ;
        RECT  24.25 6.05 24.95 6.75 ;
    END
END DFFRSX1
MACRO DFFRSX2
    CLASS CORE ;
    FOREIGN DFFRSX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 28.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  13.45 5.75 14.15 6.45 ;
        RECT  15.65 5.35 16.55 6.35 ;
        RECT  13.45 5.85 16.55 6.35 ;
        RECT  15.65 5.50 17.75 6.20 ;
        RECT  13.45 5.85 17.75 6.20 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  9.50 2.70 10.95 3.45 ;
        RECT  10.50 2.60 10.95 3.70 ;
        RECT  10.05 2.70 10.95 3.70 ;
        RECT  10.50 2.60 22.50 3.10 ;
        RECT  9.50 2.70 22.50 3.10 ;
        RECT  21.80 2.60 22.50 3.30 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  26.85 2.65 27.35 10.55 ;
        RECT  26.85 2.65 27.55 3.40 ;
        RECT  26.85 8.10 27.55 10.55 ;
        RECT  26.85 5.40 27.75 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  24.15 2.65 24.85 4.30 ;
        RECT  24.15 7.25 24.85 10.55 ;
        RECT  24.15 3.80 25.95 4.30 ;
        RECT  25.45 3.80 25.95 7.75 ;
        RECT  24.15 7.25 25.95 7.75 ;
        RECT  25.45 5.40 26.35 6.30 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.35 7.60 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.45 2.50 11.00 ;
        RECT  4.05 8.10 4.75 11.00 ;
        RECT  3.60 10.80 6.10 11.00 ;
        RECT  9.80 8.30 10.50 11.00 ;
        RECT  12.65 7.30 13.35 11.00 ;
        RECT  12.65 7.30 18.20 7.80 ;
        RECT  17.50 7.30 18.20 8.35 ;
        RECT  19.85 9.25 20.55 11.00 ;
        RECT  22.55 9.25 23.25 11.00 ;
        RECT  25.50 8.25 26.20 11.00 ;
        RECT  0.00 11.00 28.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.20 ;
        RECT  4.05 2.00 4.75 4.85 ;
        RECT  8.50 2.00 9.00 4.95 ;
        RECT  9.90 4.45 10.60 5.20 ;
        RECT  11.45 3.55 11.95 4.95 ;
        RECT  8.50 4.45 11.95 4.95 ;
        RECT  11.45 3.55 14.85 4.05 ;
        RECT  14.15 3.55 14.85 4.25 ;
        RECT  19.85 3.55 20.55 4.25 ;
        RECT  19.85 3.75 23.65 4.25 ;
        RECT  23.15 2.00 23.65 5.50 ;
        RECT  23.15 4.80 24.40 5.50 ;
        RECT  25.50 2.00 26.20 3.30 ;
        RECT  0.00 0.00 28.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.65 3.70 1.15 10.20 ;
        RECT  0.45 9.50 1.15 10.20 ;
        RECT  1.65 5.55 2.60 6.25 ;
        RECT  1.75 2.45 2.25 4.20 ;
        RECT  0.65 3.70 2.25 4.20 ;
        RECT  2.10 5.55 2.60 8.80 ;
        RECT  2.70 4.20 3.40 6.05 ;
        RECT  2.10 8.10 3.40 8.80 ;
        RECT  1.75 2.45 3.55 3.15 ;
        RECT  1.65 5.55 6.35 6.05 ;
        RECT  5.35 3.20 5.85 6.05 ;
        RECT  5.85 5.55 6.35 7.45 ;
        RECT  5.85 6.75 6.55 7.45 ;
        RECT  6.40 4.20 7.55 4.90 ;
        RECT  7.05 4.20 7.55 9.00 ;
        RECT  7.05 3.00 7.75 3.70 ;
        RECT  5.35 3.20 7.75 3.70 ;
        RECT  6.40 8.30 8.15 9.00 ;
        RECT  9.35 5.65 10.05 6.35 ;
        RECT  10.35 6.90 11.05 7.60 ;
        RECT  7.05 7.10 11.05 7.60 ;
        RECT  11.65 5.65 12.15 9.00 ;
        RECT  11.15 8.30 12.15 9.00 ;
        RECT  12.45 4.55 12.95 6.15 ;
        RECT  9.35 5.65 12.95 6.15 ;
        RECT  12.45 4.55 13.15 5.25 ;
        RECT  15.00 8.30 15.70 10.05 ;
        RECT  16.50 3.55 17.20 4.25 ;
        RECT  17.50 8.85 18.20 9.95 ;
        RECT  16.50 3.75 19.35 4.25 ;
        RECT  18.85 3.75 19.35 9.35 ;
        RECT  15.00 8.85 19.35 9.35 ;
        RECT  19.85 4.75 22.05 5.45 ;
        RECT  21.20 8.25 21.90 9.90 ;
        RECT  21.55 4.75 22.05 6.55 ;
        RECT  21.95 7.05 22.65 7.75 ;
        RECT  18.85 7.25 22.65 7.75 ;
        RECT  23.15 6.05 23.65 8.75 ;
        RECT  21.20 8.25 23.65 8.75 ;
        RECT  21.55 6.05 24.95 6.55 ;
        RECT  24.25 6.05 24.95 6.75 ;
    END
END DFFRSX2
MACRO DFFRSX4
    CLASS CORE ;
    FOREIGN DFFRSX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 30.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  13.45 5.75 14.15 6.45 ;
        RECT  15.65 5.35 16.55 6.35 ;
        RECT  13.45 5.85 16.55 6.35 ;
        RECT  15.65 5.50 17.75 6.20 ;
        RECT  13.45 5.85 17.75 6.20 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  9.50 2.70 10.95 3.45 ;
        RECT  10.50 2.60 10.95 3.70 ;
        RECT  10.05 2.70 10.95 3.70 ;
        RECT  10.50 2.60 22.50 3.10 ;
        RECT  9.50 2.70 22.50 3.10 ;
        RECT  21.80 2.60 22.50 3.30 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  28.30 2.50 29.00 4.10 ;
        RECT  28.50 2.50 29.00 10.50 ;
        RECT  28.30 5.40 29.00 10.50 ;
        RECT  28.25 5.40 29.15 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  25.60 2.50 26.10 10.50 ;
        RECT  25.60 2.50 26.30 4.10 ;
        RECT  25.60 8.10 26.30 10.50 ;
        RECT  25.45 5.40 26.35 6.30 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.35 7.60 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.45 2.50 11.00 ;
        RECT  4.05 8.10 4.75 11.00 ;
        RECT  3.60 10.80 6.10 11.00 ;
        RECT  9.80 8.30 10.50 11.00 ;
        RECT  12.65 7.30 13.35 11.00 ;
        RECT  12.65 7.30 18.20 7.80 ;
        RECT  17.50 7.30 18.20 8.35 ;
        RECT  19.85 9.25 20.55 11.00 ;
        RECT  22.55 9.25 23.25 11.00 ;
        RECT  24.25 8.10 24.95 11.00 ;
        RECT  26.95 8.10 27.65 11.00 ;
        RECT  29.65 8.10 30.35 11.00 ;
        RECT  0.00 11.00 30.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.20 ;
        RECT  4.05 2.00 4.75 4.85 ;
        RECT  8.50 2.00 9.00 4.95 ;
        RECT  9.90 4.45 10.60 5.20 ;
        RECT  11.45 3.55 11.95 4.95 ;
        RECT  8.50 4.45 11.95 4.95 ;
        RECT  11.45 3.55 14.85 4.05 ;
        RECT  14.15 3.55 14.85 4.25 ;
        RECT  19.85 3.55 20.55 4.25 ;
        RECT  24.10 2.00 24.40 5.50 ;
        RECT  23.70 3.75 24.40 5.50 ;
        RECT  24.10 2.00 24.80 4.25 ;
        RECT  19.85 3.75 24.80 4.25 ;
        RECT  26.95 2.00 27.65 4.10 ;
        RECT  29.65 2.00 30.35 4.10 ;
        RECT  0.00 0.00 30.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.65 3.70 1.15 10.20 ;
        RECT  0.45 9.50 1.15 10.20 ;
        RECT  1.65 5.55 2.60 6.25 ;
        RECT  1.75 2.45 2.25 4.20 ;
        RECT  0.65 3.70 2.25 4.20 ;
        RECT  2.10 5.55 2.60 8.80 ;
        RECT  2.70 4.20 3.40 6.05 ;
        RECT  2.10 8.10 3.40 8.80 ;
        RECT  1.75 2.45 3.55 3.15 ;
        RECT  1.65 5.55 6.35 6.05 ;
        RECT  5.35 3.20 5.85 6.05 ;
        RECT  5.85 5.55 6.35 7.45 ;
        RECT  5.85 6.75 6.55 7.45 ;
        RECT  6.40 4.20 7.55 4.90 ;
        RECT  7.05 4.20 7.55 9.00 ;
        RECT  7.05 3.00 7.75 3.70 ;
        RECT  5.35 3.20 7.75 3.70 ;
        RECT  6.40 8.30 8.15 9.00 ;
        RECT  9.35 5.65 10.05 6.35 ;
        RECT  10.35 6.90 11.05 7.60 ;
        RECT  7.05 7.10 11.05 7.60 ;
        RECT  11.65 5.65 12.15 9.00 ;
        RECT  11.15 8.30 12.15 9.00 ;
        RECT  12.45 4.55 12.95 6.15 ;
        RECT  9.35 5.65 12.95 6.15 ;
        RECT  12.45 4.55 13.15 5.25 ;
        RECT  15.00 8.30 15.70 10.05 ;
        RECT  16.50 3.55 17.20 4.25 ;
        RECT  17.50 8.85 18.20 9.95 ;
        RECT  16.50 3.75 19.35 4.25 ;
        RECT  18.85 3.75 19.35 9.35 ;
        RECT  15.00 8.85 19.35 9.35 ;
        RECT  19.85 4.75 22.05 5.45 ;
        RECT  21.20 8.25 21.90 9.90 ;
        RECT  21.55 4.75 22.05 6.55 ;
        RECT  21.95 7.05 22.65 7.75 ;
        RECT  18.85 7.25 22.65 7.75 ;
        RECT  23.15 6.05 23.65 8.75 ;
        RECT  21.20 8.25 23.65 8.75 ;
        RECT  21.55 6.05 24.95 6.55 ;
        RECT  24.25 6.05 24.95 6.75 ;
    END
END DFFRSX4
MACRO DFFRX1
    CLASS CORE ;
    FOREIGN DFFRX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 25.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  9.15 2.45 9.85 3.45 ;
        RECT  15.65 2.45 16.55 3.75 ;
        RECT  9.15 2.45 18.60 2.95 ;
        RECT  17.90 2.45 18.60 3.15 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  24.05 3.75 24.55 9.50 ;
        RECT  24.05 3.75 24.75 6.30 ;
        RECT  24.05 7.85 24.75 9.50 ;
        RECT  24.05 5.40 24.95 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  21.35 3.75 22.05 5.40 ;
        RECT  21.35 7.00 22.05 9.50 ;
        RECT  21.35 4.90 23.15 5.40 ;
        RECT  22.65 4.90 23.15 7.50 ;
        RECT  21.35 7.00 23.15 7.50 ;
        RECT  22.65 5.40 23.55 6.30 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.35 7.60 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.50 2.50 11.00 ;
        RECT  4.05 8.10 4.75 11.00 ;
        RECT  3.60 10.80 6.10 11.00 ;
        RECT  9.80 8.30 10.50 11.00 ;
        RECT  12.30 9.70 13.00 11.00 ;
        RECT  17.15 9.30 17.85 11.00 ;
        RECT  19.85 9.30 20.55 11.00 ;
        RECT  22.70 8.00 23.40 11.00 ;
        RECT  0.00 11.00 25.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.20 ;
        RECT  4.05 2.00 4.75 4.85 ;
        RECT  8.20 2.00 8.70 4.40 ;
        RECT  8.20 3.90 10.80 4.40 ;
        RECT  10.30 3.60 10.80 5.20 ;
        RECT  9.90 3.90 10.80 5.20 ;
        RECT  10.30 3.60 13.45 4.10 ;
        RECT  8.20 3.90 13.45 4.10 ;
        RECT  12.75 3.60 13.45 5.20 ;
        RECT  17.60 3.60 18.15 5.20 ;
        RECT  17.45 4.45 18.15 5.20 ;
        RECT  19.05 2.00 19.55 4.10 ;
        RECT  17.60 3.60 19.55 4.10 ;
        RECT  22.70 2.00 23.40 4.40 ;
        RECT  0.00 0.00 25.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.65 3.70 1.15 10.20 ;
        RECT  0.45 9.50 1.15 10.20 ;
        RECT  1.65 5.55 2.60 6.25 ;
        RECT  1.75 2.45 2.25 4.20 ;
        RECT  0.65 3.70 2.25 4.20 ;
        RECT  2.10 5.55 2.60 8.75 ;
        RECT  2.70 4.20 3.40 6.05 ;
        RECT  2.10 8.05 3.40 8.75 ;
        RECT  1.75 2.45 3.55 3.15 ;
        RECT  1.65 5.55 6.35 6.05 ;
        RECT  5.35 3.20 5.85 6.05 ;
        RECT  5.85 5.55 6.35 7.45 ;
        RECT  5.85 6.75 6.55 7.45 ;
        RECT  6.40 4.20 7.55 4.90 ;
        RECT  7.05 4.20 7.55 9.00 ;
        RECT  7.05 3.00 7.75 3.70 ;
        RECT  5.35 3.20 7.75 3.70 ;
        RECT  6.40 8.30 8.15 9.00 ;
        RECT  9.35 5.65 10.05 6.35 ;
        RECT  10.25 6.90 10.95 7.60 ;
        RECT  7.05 7.10 10.95 7.60 ;
        RECT  11.25 4.55 11.95 6.15 ;
        RECT  9.35 5.65 11.95 6.15 ;
        RECT  11.45 4.55 11.95 9.00 ;
        RECT  11.15 8.25 11.95 9.00 ;
        RECT  15.10 4.50 15.50 10.05 ;
        RECT  14.80 7.30 15.50 10.05 ;
        RECT  15.10 4.50 15.60 7.90 ;
        RECT  15.10 4.50 15.80 5.20 ;
        RECT  16.80 5.75 17.50 6.45 ;
        RECT  18.50 8.35 19.20 9.95 ;
        RECT  18.90 7.20 19.60 7.90 ;
        RECT  14.80 7.30 19.60 7.90 ;
        RECT  16.80 5.75 20.55 6.25 ;
        RECT  19.85 4.55 20.55 6.25 ;
        RECT  16.80 5.85 22.15 6.25 ;
        RECT  20.05 4.55 20.55 8.85 ;
        RECT  18.50 8.35 20.55 8.85 ;
        RECT  20.05 5.85 22.15 6.55 ;
    END
END DFFRX1
MACRO DFFRX2
    CLASS CORE ;
    FOREIGN DFFRX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 25.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  9.15 2.45 9.85 3.45 ;
        RECT  15.65 2.45 16.55 3.75 ;
        RECT  9.15 2.45 18.60 2.95 ;
        RECT  17.90 2.45 18.60 3.15 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  24.05 2.70 24.55 10.55 ;
        RECT  24.05 2.70 24.75 6.30 ;
        RECT  24.05 7.85 24.75 10.55 ;
        RECT  24.05 5.40 24.95 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  21.35 2.70 22.05 5.40 ;
        RECT  21.35 7.00 22.05 10.55 ;
        RECT  21.35 4.90 23.15 5.40 ;
        RECT  22.65 4.90 23.15 7.50 ;
        RECT  21.35 7.00 23.15 7.50 ;
        RECT  22.65 5.40 23.55 6.30 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.35 7.60 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.45 2.50 11.00 ;
        RECT  4.05 8.05 4.75 11.00 ;
        RECT  3.60 10.95 6.10 11.00 ;
        RECT  9.80 8.30 10.50 11.00 ;
        RECT  12.30 9.70 13.00 11.00 ;
        RECT  17.15 9.30 17.85 11.00 ;
        RECT  19.85 9.30 20.55 11.00 ;
        RECT  22.70 8.00 23.40 11.00 ;
        RECT  0.00 11.00 25.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.20 ;
        RECT  4.05 2.00 4.75 4.85 ;
        RECT  8.20 2.00 8.70 4.40 ;
        RECT  8.20 3.90 10.80 4.40 ;
        RECT  10.30 3.60 10.80 5.20 ;
        RECT  9.90 3.90 10.80 5.20 ;
        RECT  10.30 3.60 13.45 4.10 ;
        RECT  8.20 3.90 13.45 4.10 ;
        RECT  12.75 3.60 13.45 5.20 ;
        RECT  17.60 3.60 18.15 5.20 ;
        RECT  17.45 4.45 18.15 5.20 ;
        RECT  19.05 2.00 19.55 4.10 ;
        RECT  17.60 3.60 19.55 4.10 ;
        RECT  22.70 2.00 23.40 4.40 ;
        RECT  0.00 0.00 25.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.65 3.70 1.15 10.15 ;
        RECT  0.45 9.45 1.15 10.15 ;
        RECT  1.65 5.55 2.60 6.25 ;
        RECT  1.75 2.45 2.25 4.20 ;
        RECT  0.65 3.70 2.25 4.20 ;
        RECT  2.10 5.55 2.60 8.75 ;
        RECT  2.70 4.20 3.40 6.05 ;
        RECT  2.10 8.05 3.40 8.75 ;
        RECT  1.75 2.45 3.55 3.15 ;
        RECT  1.65 5.55 6.35 6.05 ;
        RECT  5.35 3.20 5.85 6.05 ;
        RECT  5.85 5.55 6.35 7.45 ;
        RECT  5.85 6.75 6.55 7.45 ;
        RECT  6.40 4.20 7.55 4.90 ;
        RECT  7.05 4.20 7.55 9.00 ;
        RECT  7.05 3.00 7.75 3.70 ;
        RECT  5.35 3.20 7.75 3.70 ;
        RECT  6.40 8.30 8.15 9.00 ;
        RECT  9.35 5.65 10.05 6.35 ;
        RECT  10.25 6.90 10.95 7.60 ;
        RECT  7.05 7.10 10.95 7.60 ;
        RECT  11.25 4.55 11.95 6.15 ;
        RECT  9.35 5.65 11.95 6.15 ;
        RECT  11.45 4.55 11.95 9.00 ;
        RECT  11.15 8.25 11.95 9.00 ;
        RECT  15.10 4.50 15.50 10.05 ;
        RECT  14.80 7.30 15.50 10.05 ;
        RECT  15.10 4.50 15.60 7.90 ;
        RECT  15.10 4.50 15.80 5.20 ;
        RECT  16.80 5.75 17.50 6.45 ;
        RECT  18.50 8.35 19.20 9.95 ;
        RECT  18.90 7.20 19.60 7.90 ;
        RECT  14.80 7.30 19.60 7.90 ;
        RECT  16.80 5.75 20.55 6.25 ;
        RECT  19.85 4.55 20.55 6.25 ;
        RECT  16.80 5.85 22.15 6.25 ;
        RECT  20.05 4.55 20.55 8.85 ;
        RECT  18.50 8.35 20.55 8.85 ;
        RECT  20.05 5.85 22.15 6.55 ;
    END
END DFFRX2
MACRO DFFRX4
    CLASS CORE ;
    FOREIGN DFFRX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 28.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  9.15 2.45 9.85 3.45 ;
        RECT  15.65 2.45 16.55 3.75 ;
        RECT  9.15 2.45 18.60 2.95 ;
        RECT  17.90 2.45 18.60 3.15 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  25.50 2.90 26.20 10.55 ;
        RECT  25.45 5.40 26.35 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  22.80 2.90 23.50 10.55 ;
        RECT  22.65 5.40 23.55 6.30 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.55 5.35 7.60 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.55 3.95 7.60 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.35 2.50 11.00 ;
        RECT  4.05 8.05 4.75 11.00 ;
        RECT  3.60 10.75 6.10 11.00 ;
        RECT  9.80 8.30 10.50 11.00 ;
        RECT  12.30 9.70 13.00 11.00 ;
        RECT  17.15 9.30 17.85 11.00 ;
        RECT  19.85 9.30 20.55 11.00 ;
        RECT  21.45 7.85 22.15 11.00 ;
        RECT  24.15 7.85 24.85 11.00 ;
        RECT  26.85 7.85 27.55 11.00 ;
        RECT  0.00 11.00 28.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.20 ;
        RECT  4.05 2.00 4.75 4.85 ;
        RECT  8.20 2.00 8.70 4.40 ;
        RECT  8.20 3.90 10.80 4.40 ;
        RECT  10.30 3.60 10.80 5.20 ;
        RECT  9.90 3.90 10.80 5.20 ;
        RECT  10.30 3.60 13.45 4.10 ;
        RECT  8.20 3.90 13.45 4.10 ;
        RECT  12.75 3.60 13.45 5.20 ;
        RECT  17.60 3.60 18.15 5.20 ;
        RECT  17.45 4.45 18.15 5.20 ;
        RECT  19.05 2.00 19.55 4.10 ;
        RECT  17.60 3.60 19.55 4.10 ;
        RECT  21.45 2.00 22.15 4.50 ;
        RECT  24.15 2.00 24.85 4.50 ;
        RECT  26.85 2.00 27.55 4.50 ;
        RECT  0.00 0.00 28.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.65 3.70 1.15 10.15 ;
        RECT  0.45 9.45 1.15 10.15 ;
        RECT  1.65 5.55 2.60 6.25 ;
        RECT  1.75 2.45 2.25 4.20 ;
        RECT  0.65 3.70 2.25 4.20 ;
        RECT  2.10 5.55 2.60 8.75 ;
        RECT  2.70 4.20 3.40 6.05 ;
        RECT  2.10 8.05 3.40 8.75 ;
        RECT  1.75 2.45 3.55 3.15 ;
        RECT  1.65 5.55 6.35 6.05 ;
        RECT  5.35 3.20 5.85 6.05 ;
        RECT  5.85 5.55 6.35 7.45 ;
        RECT  5.85 6.75 6.55 7.45 ;
        RECT  6.40 4.20 7.55 4.90 ;
        RECT  7.05 4.20 7.55 9.00 ;
        RECT  7.05 3.00 7.75 3.70 ;
        RECT  5.35 3.20 7.75 3.70 ;
        RECT  6.40 8.30 8.15 9.00 ;
        RECT  9.35 5.65 10.05 6.35 ;
        RECT  10.25 6.90 10.95 7.60 ;
        RECT  7.05 7.10 10.95 7.60 ;
        RECT  11.25 4.55 11.95 6.15 ;
        RECT  9.35 5.65 11.95 6.15 ;
        RECT  11.45 4.55 11.95 9.00 ;
        RECT  11.15 8.25 11.95 9.00 ;
        RECT  15.10 4.50 15.50 10.05 ;
        RECT  14.80 7.30 15.50 10.05 ;
        RECT  15.10 4.50 15.60 7.90 ;
        RECT  15.10 4.50 15.80 5.20 ;
        RECT  16.80 5.75 17.50 6.45 ;
        RECT  18.50 8.35 19.20 9.95 ;
        RECT  18.90 7.20 19.60 7.90 ;
        RECT  14.80 7.30 19.60 7.90 ;
        RECT  16.80 5.75 20.55 6.25 ;
        RECT  19.85 4.55 20.55 6.25 ;
        RECT  16.80 6.00 22.15 6.25 ;
        RECT  20.05 4.55 20.55 8.85 ;
        RECT  18.50 8.35 20.55 8.85 ;
        RECT  20.05 6.00 22.15 6.50 ;
        RECT  21.45 6.00 22.15 6.70 ;
    END
END DFFRX4
MACRO DFFSX1
    CLASS CORE ;
    FOREIGN DFFSX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  11.45 7.05 12.15 8.40 ;
        RECT  12.85 6.70 13.75 7.60 ;
        RECT  13.25 5.45 13.75 7.60 ;
        RECT  11.45 7.05 13.75 7.60 ;
        RECT  13.90 5.25 14.60 5.95 ;
        RECT  13.25 5.45 14.60 5.95 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  19.95 3.75 20.65 4.45 ;
        RECT  20.10 3.75 20.65 8.85 ;
        RECT  19.95 7.15 20.65 8.85 ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  22.65 3.75 23.35 4.45 ;
        RECT  22.85 3.75 23.35 8.85 ;
        RECT  22.65 7.15 23.35 8.85 ;
        RECT  22.65 5.40 23.55 6.30 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.35 7.60 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.45 2.50 11.00 ;
        RECT  4.05 8.05 4.75 11.00 ;
        RECT  3.30 10.75 6.95 11.00 ;
        RECT  8.75 8.00 9.45 11.00 ;
        RECT  8.00 10.65 9.60 11.00 ;
        RECT  12.05 8.90 12.75 11.00 ;
        RECT  17.05 7.40 17.75 11.00 ;
        RECT  21.30 7.15 22.00 11.00 ;
        RECT  17.05 10.70 23.35 11.00 ;
        RECT  0.00 11.00 23.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.20 ;
        RECT  4.05 2.00 4.75 4.90 ;
        RECT  8.15 2.00 9.75 3.30 ;
        RECT  9.05 2.00 9.75 4.90 ;
        RECT  11.20 2.00 11.90 3.25 ;
        RECT  17.05 2.00 17.75 3.95 ;
        RECT  21.30 2.00 22.00 4.45 ;
        RECT  0.00 0.00 23.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.65 3.70 1.15 10.15 ;
        RECT  0.45 9.45 1.15 10.15 ;
        RECT  1.65 5.55 2.60 6.25 ;
        RECT  1.75 2.45 2.25 4.20 ;
        RECT  0.65 3.70 2.25 4.20 ;
        RECT  2.10 5.55 2.60 8.75 ;
        RECT  2.70 4.20 3.40 6.05 ;
        RECT  2.10 8.05 3.40 8.75 ;
        RECT  1.75 2.45 3.55 3.15 ;
        RECT  1.65 5.55 6.35 6.05 ;
        RECT  5.35 3.20 5.85 6.05 ;
        RECT  5.85 5.55 6.35 7.50 ;
        RECT  5.85 6.80 6.55 7.50 ;
        RECT  6.40 4.20 7.50 4.90 ;
        RECT  7.00 4.20 7.10 9.65 ;
        RECT  6.40 8.05 7.10 9.65 ;
        RECT  7.00 4.20 7.50 8.75 ;
        RECT  6.40 8.05 7.50 8.75 ;
        RECT  7.00 3.00 7.70 3.70 ;
        RECT  5.35 3.20 7.70 3.70 ;
        RECT  8.30 5.45 9.00 6.15 ;
        RECT  7.00 6.70 9.95 7.20 ;
        RECT  9.25 6.70 9.95 7.40 ;
        RECT  8.30 5.45 10.95 5.95 ;
        RECT  10.45 4.45 10.95 9.70 ;
        RECT  10.45 9.00 11.25 9.70 ;
        RECT  11.55 4.25 12.25 4.95 ;
        RECT  10.45 4.45 12.25 4.95 ;
        RECT  13.70 3.30 14.40 4.00 ;
        RECT  13.70 3.45 15.60 4.00 ;
        RECT  14.55 7.20 15.10 10.50 ;
        RECT  14.40 8.75 15.10 10.50 ;
        RECT  15.10 3.45 15.60 7.90 ;
        RECT  14.55 7.20 15.60 7.90 ;
        RECT  16.60 4.45 17.30 5.15 ;
        RECT  17.40 5.70 18.10 6.40 ;
        RECT  15.10 5.90 18.10 6.40 ;
        RECT  18.40 3.25 19.10 3.95 ;
        RECT  16.60 4.45 19.10 4.95 ;
        RECT  18.60 3.25 19.10 10.10 ;
        RECT  18.40 7.40 19.10 10.10 ;
    END
END DFFSX1
MACRO DFFSX2
    CLASS CORE ;
    FOREIGN DFFSX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  11.45 7.05 12.15 8.40 ;
        RECT  12.85 6.70 13.75 7.60 ;
        RECT  13.25 5.45 13.75 7.60 ;
        RECT  11.45 7.05 13.75 7.60 ;
        RECT  13.90 5.25 14.60 5.95 ;
        RECT  13.25 5.45 14.60 5.95 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  19.95 2.70 20.65 4.50 ;
        RECT  20.10 2.70 20.65 10.55 ;
        RECT  19.95 7.10 20.65 10.55 ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  22.65 2.70 23.35 4.50 ;
        RECT  22.85 2.70 23.35 10.55 ;
        RECT  22.65 7.10 23.35 10.55 ;
        RECT  22.65 5.40 23.55 6.30 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.35 7.60 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.45 2.50 11.00 ;
        RECT  4.05 8.05 4.75 11.00 ;
        RECT  3.30 10.75 6.95 11.00 ;
        RECT  8.75 7.95 9.45 11.00 ;
        RECT  8.00 10.65 9.60 11.00 ;
        RECT  12.05 8.90 12.75 11.00 ;
        RECT  17.05 7.40 17.75 11.00 ;
        RECT  21.30 7.10 22.00 11.00 ;
        RECT  0.00 11.00 23.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.20 ;
        RECT  4.05 2.00 4.75 4.90 ;
        RECT  8.15 2.00 9.75 3.30 ;
        RECT  9.05 2.00 9.75 4.90 ;
        RECT  11.20 2.00 11.90 3.25 ;
        RECT  17.05 2.00 17.75 3.95 ;
        RECT  21.30 2.00 22.00 4.50 ;
        RECT  0.00 0.00 23.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.65 3.70 1.15 10.15 ;
        RECT  0.45 9.45 1.15 10.15 ;
        RECT  1.65 5.55 2.60 6.25 ;
        RECT  1.75 2.45 2.25 4.20 ;
        RECT  0.65 3.70 2.25 4.20 ;
        RECT  2.10 5.55 2.60 8.75 ;
        RECT  2.70 4.20 3.40 6.05 ;
        RECT  2.10 8.05 3.40 8.75 ;
        RECT  1.75 2.45 3.55 3.15 ;
        RECT  1.65 5.55 6.35 6.05 ;
        RECT  5.35 3.20 5.85 6.05 ;
        RECT  5.85 5.55 6.35 7.50 ;
        RECT  5.85 6.80 6.55 7.50 ;
        RECT  6.40 4.20 7.50 4.90 ;
        RECT  7.00 4.20 7.10 9.75 ;
        RECT  6.40 8.05 7.10 9.75 ;
        RECT  7.00 4.20 7.50 8.85 ;
        RECT  6.40 8.05 7.50 8.85 ;
        RECT  7.00 3.00 7.70 3.70 ;
        RECT  5.35 3.20 7.70 3.70 ;
        RECT  8.30 5.45 9.00 6.15 ;
        RECT  7.00 6.70 9.95 7.20 ;
        RECT  9.25 6.70 9.95 7.40 ;
        RECT  8.30 5.45 10.95 5.95 ;
        RECT  10.45 4.45 10.95 9.70 ;
        RECT  10.45 9.00 11.25 9.70 ;
        RECT  11.55 4.25 12.25 4.95 ;
        RECT  10.45 4.45 12.25 4.95 ;
        RECT  13.70 3.30 14.40 4.00 ;
        RECT  13.70 3.45 15.60 4.00 ;
        RECT  14.55 7.20 15.10 10.50 ;
        RECT  14.40 8.75 15.10 10.50 ;
        RECT  15.10 3.45 15.60 7.90 ;
        RECT  14.55 7.20 15.60 7.90 ;
        RECT  16.60 4.45 17.30 5.15 ;
        RECT  17.40 5.70 18.10 6.40 ;
        RECT  15.10 5.90 18.10 6.40 ;
        RECT  18.40 3.25 19.10 3.95 ;
        RECT  16.60 4.45 19.10 4.95 ;
        RECT  18.60 3.25 19.10 10.55 ;
        RECT  18.40 7.40 19.10 10.55 ;
    END
END DFFSX2
MACRO DFFSX4
    CLASS CORE ;
    FOREIGN DFFSX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 26.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  11.45 7.05 12.15 8.40 ;
        RECT  12.85 6.70 13.75 7.60 ;
        RECT  13.25 5.45 13.75 7.60 ;
        RECT  11.45 7.05 13.75 7.60 ;
        RECT  13.90 5.25 14.60 5.95 ;
        RECT  13.25 5.45 14.60 5.95 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  21.40 2.70 22.10 10.50 ;
        RECT  21.25 5.40 22.15 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  24.10 2.70 24.80 10.50 ;
        RECT  24.05 5.40 24.95 6.30 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.35 7.60 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.45 2.50 11.00 ;
        RECT  4.05 8.05 4.75 11.00 ;
        RECT  3.30 10.75 6.95 11.00 ;
        RECT  8.75 8.00 9.45 11.00 ;
        RECT  8.00 10.65 9.60 11.00 ;
        RECT  12.05 8.90 12.75 11.00 ;
        RECT  17.05 7.40 17.75 11.00 ;
        RECT  20.05 7.10 20.75 11.00 ;
        RECT  22.75 7.10 23.45 11.00 ;
        RECT  25.45 7.10 26.15 11.00 ;
        RECT  0.00 11.00 26.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.20 ;
        RECT  4.05 2.00 4.75 4.90 ;
        RECT  8.15 2.00 9.75 3.30 ;
        RECT  9.05 2.00 9.75 4.90 ;
        RECT  11.20 2.00 11.90 3.25 ;
        RECT  17.05 2.00 17.75 3.95 ;
        RECT  20.05 2.00 20.75 4.50 ;
        RECT  22.75 2.00 23.45 4.50 ;
        RECT  25.45 2.00 26.15 4.50 ;
        RECT  0.00 0.00 26.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.65 3.70 1.15 10.15 ;
        RECT  0.45 9.35 1.15 10.15 ;
        RECT  1.65 5.55 2.60 6.25 ;
        RECT  1.75 2.45 2.25 4.20 ;
        RECT  0.65 3.70 2.25 4.20 ;
        RECT  2.10 5.55 2.60 8.75 ;
        RECT  2.70 4.20 3.40 6.05 ;
        RECT  2.10 8.05 3.40 8.75 ;
        RECT  1.75 2.45 3.55 3.15 ;
        RECT  1.65 5.55 6.35 6.05 ;
        RECT  5.35 3.20 5.85 6.05 ;
        RECT  5.85 5.55 6.35 7.50 ;
        RECT  5.85 6.80 6.55 7.50 ;
        RECT  6.40 4.20 7.50 4.90 ;
        RECT  7.00 4.20 7.10 9.70 ;
        RECT  6.40 8.05 7.10 9.70 ;
        RECT  7.00 4.20 7.50 8.75 ;
        RECT  6.40 8.05 7.50 8.75 ;
        RECT  7.00 3.00 7.70 3.70 ;
        RECT  5.35 3.20 7.70 3.70 ;
        RECT  8.30 5.45 9.00 6.15 ;
        RECT  7.00 6.70 9.95 7.20 ;
        RECT  9.25 6.70 9.95 7.40 ;
        RECT  8.30 5.45 10.95 5.95 ;
        RECT  10.45 4.45 10.95 9.70 ;
        RECT  10.45 9.00 11.25 9.70 ;
        RECT  11.55 4.25 12.25 4.95 ;
        RECT  10.45 4.45 12.25 4.95 ;
        RECT  13.70 3.30 14.40 4.00 ;
        RECT  13.70 3.45 15.60 4.00 ;
        RECT  14.55 7.20 15.10 10.50 ;
        RECT  14.40 8.75 15.10 10.50 ;
        RECT  15.10 3.45 15.60 7.90 ;
        RECT  14.55 7.20 15.60 7.90 ;
        RECT  16.60 4.45 17.30 5.15 ;
        RECT  17.40 5.70 18.10 6.40 ;
        RECT  15.10 5.90 18.10 6.40 ;
        RECT  18.40 3.25 19.10 4.95 ;
        RECT  16.60 4.45 19.60 4.95 ;
        RECT  18.60 3.25 19.10 10.55 ;
        RECT  18.40 7.40 19.10 10.55 ;
        RECT  18.60 4.45 19.60 5.15 ;
    END
END DFFSX4
MACRO DFFX1
    CLASS CORE ;
    FOREIGN DFFX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  17.15 3.75 17.85 4.45 ;
        RECT  17.30 3.75 17.85 8.85 ;
        RECT  17.15 7.15 17.85 8.85 ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  19.85 3.75 20.55 4.45 ;
        RECT  20.05 3.75 20.55 8.85 ;
        RECT  19.85 7.15 20.55 8.85 ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.35 7.60 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.45 2.50 11.00 ;
        RECT  4.05 8.05 4.75 11.00 ;
        RECT  3.30 10.70 6.95 11.00 ;
        RECT  8.75 7.90 9.45 11.00 ;
        RECT  8.00 10.50 10.15 11.00 ;
        RECT  10.95 10.40 11.65 11.00 ;
        RECT  14.25 7.40 14.95 8.15 ;
        RECT  14.45 7.40 14.95 11.00 ;
        RECT  14.45 10.15 16.50 11.00 ;
        RECT  18.50 7.15 19.20 11.00 ;
        RECT  17.30 10.70 20.55 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.20 ;
        RECT  4.05 2.00 4.75 4.85 ;
        RECT  8.75 2.00 9.45 4.85 ;
        RECT  8.75 2.00 10.05 3.15 ;
        RECT  14.25 2.00 14.95 3.95 ;
        RECT  18.50 2.00 19.20 4.45 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.65 3.70 1.15 10.15 ;
        RECT  0.45 9.45 1.15 10.15 ;
        RECT  1.65 5.55 2.60 6.25 ;
        RECT  1.75 2.45 2.25 4.20 ;
        RECT  0.65 3.70 2.25 4.20 ;
        RECT  2.10 5.55 2.60 8.75 ;
        RECT  2.70 4.10 3.40 6.15 ;
        RECT  1.65 5.55 3.40 6.15 ;
        RECT  2.10 8.05 3.40 8.75 ;
        RECT  1.75 2.45 3.55 3.15 ;
        RECT  1.65 5.65 6.30 6.15 ;
        RECT  5.80 3.15 5.85 7.45 ;
        RECT  5.35 3.15 5.85 6.15 ;
        RECT  5.80 5.65 6.30 7.45 ;
        RECT  5.80 6.75 6.50 7.45 ;
        RECT  6.40 4.15 7.50 4.85 ;
        RECT  7.00 4.15 7.10 9.75 ;
        RECT  6.40 8.00 7.10 9.75 ;
        RECT  7.00 4.15 7.50 8.50 ;
        RECT  6.40 8.00 7.50 8.50 ;
        RECT  7.00 2.95 7.70 3.65 ;
        RECT  5.35 3.15 7.70 3.65 ;
        RECT  8.30 5.45 9.00 6.15 ;
        RECT  7.00 6.75 9.95 7.25 ;
        RECT  9.25 6.75 9.95 7.45 ;
        RECT  8.30 5.45 10.95 5.95 ;
        RECT  10.45 4.15 10.80 8.60 ;
        RECT  10.10 4.15 10.80 5.95 ;
        RECT  10.45 5.45 10.95 8.60 ;
        RECT  10.25 7.90 10.95 8.60 ;
        RECT  11.90 3.30 12.60 4.00 ;
        RECT  12.10 3.30 12.60 10.15 ;
        RECT  12.10 9.65 14.00 10.15 ;
        RECT  13.30 9.65 14.00 10.35 ;
        RECT  13.80 4.45 14.50 5.15 ;
        RECT  14.60 5.70 15.30 6.40 ;
        RECT  12.10 5.90 15.30 6.40 ;
        RECT  15.60 3.25 16.30 3.95 ;
        RECT  13.80 4.45 16.30 4.95 ;
        RECT  15.60 7.40 16.30 8.15 ;
        RECT  15.80 3.25 16.30 9.65 ;
        RECT  15.80 8.95 16.65 9.65 ;
    END
END DFFX1
MACRO DFFX2
    CLASS CORE ;
    FOREIGN DFFX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  17.15 2.70 17.85 4.45 ;
        RECT  17.30 2.70 17.85 9.60 ;
        RECT  17.15 7.10 17.85 9.60 ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  19.85 2.70 20.55 4.45 ;
        RECT  20.05 2.70 20.55 10.50 ;
        RECT  19.85 7.10 20.55 10.50 ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.35 7.60 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.45 2.50 11.00 ;
        RECT  4.05 8.05 4.75 11.00 ;
        RECT  3.30 10.60 6.95 11.00 ;
        RECT  8.75 7.90 9.45 11.00 ;
        RECT  8.00 10.50 10.15 11.00 ;
        RECT  10.95 10.40 11.65 11.00 ;
        RECT  14.25 7.10 14.95 7.85 ;
        RECT  14.45 7.10 14.95 11.00 ;
        RECT  14.45 10.20 16.50 11.00 ;
        RECT  18.50 7.10 19.20 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.20 ;
        RECT  4.05 2.00 4.75 4.85 ;
        RECT  8.80 2.00 9.50 4.85 ;
        RECT  8.80 2.00 10.10 3.10 ;
        RECT  14.25 2.00 14.95 3.95 ;
        RECT  18.50 2.00 19.20 4.45 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.65 3.70 1.15 10.15 ;
        RECT  0.45 9.45 1.15 10.15 ;
        RECT  1.65 5.55 2.60 6.25 ;
        RECT  1.75 2.45 2.25 4.20 ;
        RECT  0.65 3.70 2.25 4.20 ;
        RECT  2.10 5.55 2.60 8.75 ;
        RECT  2.70 4.15 3.40 6.05 ;
        RECT  2.10 8.05 3.40 8.75 ;
        RECT  1.75 2.45 3.55 3.15 ;
        RECT  1.65 5.55 6.30 6.05 ;
        RECT  5.80 3.15 5.85 7.45 ;
        RECT  5.35 3.15 5.85 6.05 ;
        RECT  5.80 5.55 6.30 7.45 ;
        RECT  5.80 6.75 6.50 7.45 ;
        RECT  6.40 4.15 7.50 4.85 ;
        RECT  7.00 4.15 7.10 9.60 ;
        RECT  6.40 8.00 7.10 9.60 ;
        RECT  7.00 4.15 7.50 8.50 ;
        RECT  6.40 8.00 7.50 8.50 ;
        RECT  7.00 2.95 7.70 3.65 ;
        RECT  5.35 3.15 7.70 3.65 ;
        RECT  8.30 5.45 9.00 6.15 ;
        RECT  7.00 6.75 9.95 7.25 ;
        RECT  9.25 6.75 9.95 7.45 ;
        RECT  10.25 4.15 10.95 4.85 ;
        RECT  8.30 5.45 10.95 5.95 ;
        RECT  10.45 4.15 10.95 8.60 ;
        RECT  10.25 7.90 10.95 8.60 ;
        RECT  11.90 3.30 12.60 4.00 ;
        RECT  12.10 3.30 12.60 10.15 ;
        RECT  12.10 9.65 14.00 10.15 ;
        RECT  13.30 9.65 14.00 10.35 ;
        RECT  13.80 4.45 14.50 5.15 ;
        RECT  14.60 5.70 15.30 6.40 ;
        RECT  12.10 5.90 15.30 6.40 ;
        RECT  15.60 3.25 16.30 3.95 ;
        RECT  13.80 4.45 16.30 4.95 ;
        RECT  15.60 7.40 16.30 8.15 ;
        RECT  15.80 3.25 16.30 9.65 ;
        RECT  15.80 8.95 16.65 9.65 ;
    END
END DFFX2
MACRO DFFX4
    CLASS CORE ;
    FOREIGN DFFX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  18.60 2.70 19.30 10.50 ;
        RECT  18.45 5.40 19.35 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  21.30 2.70 22.00 10.50 ;
        RECT  21.25 5.40 22.15 6.30 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.35 7.60 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.45 2.50 11.00 ;
        RECT  4.05 8.05 4.75 11.00 ;
        RECT  3.30 10.70 6.95 11.00 ;
        RECT  8.75 7.90 9.45 11.00 ;
        RECT  8.00 10.50 10.15 11.00 ;
        RECT  10.95 10.40 11.65 11.00 ;
        RECT  14.25 7.10 14.95 7.85 ;
        RECT  14.45 7.10 14.95 11.00 ;
        RECT  17.25 7.10 17.95 11.00 ;
        RECT  19.95 7.10 20.65 11.00 ;
        RECT  22.65 7.10 23.35 11.00 ;
        RECT  0.00 11.00 23.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.20 ;
        RECT  4.05 2.00 4.75 4.85 ;
        RECT  8.80 2.00 9.50 4.85 ;
        RECT  8.80 2.00 10.10 3.15 ;
        RECT  14.25 2.00 14.95 3.95 ;
        RECT  17.25 2.00 17.95 4.50 ;
        RECT  19.95 2.00 20.65 4.50 ;
        RECT  22.65 2.00 23.35 4.50 ;
        RECT  0.00 0.00 23.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.65 3.70 1.15 10.25 ;
        RECT  0.45 9.45 1.15 10.25 ;
        RECT  1.65 5.55 2.60 6.25 ;
        RECT  1.75 2.45 2.25 4.20 ;
        RECT  0.65 3.70 2.25 4.20 ;
        RECT  2.10 5.55 2.60 8.75 ;
        RECT  2.70 4.15 3.40 6.05 ;
        RECT  2.10 8.05 3.40 8.75 ;
        RECT  1.75 2.45 3.55 3.15 ;
        RECT  1.65 5.55 6.30 6.05 ;
        RECT  5.80 3.15 5.85 7.45 ;
        RECT  5.35 3.15 5.85 6.05 ;
        RECT  5.80 5.55 6.30 7.45 ;
        RECT  5.80 6.75 6.50 7.45 ;
        RECT  6.40 4.15 7.50 4.85 ;
        RECT  7.00 4.15 7.10 9.60 ;
        RECT  6.40 8.00 7.10 9.60 ;
        RECT  7.00 4.15 7.50 8.50 ;
        RECT  6.40 8.00 7.50 8.50 ;
        RECT  7.00 2.95 7.70 3.65 ;
        RECT  5.35 3.15 7.70 3.65 ;
        RECT  8.30 5.45 9.00 6.15 ;
        RECT  7.00 6.75 9.95 7.25 ;
        RECT  9.25 6.75 9.95 7.45 ;
        RECT  10.25 4.15 10.95 4.85 ;
        RECT  8.30 5.45 10.95 5.95 ;
        RECT  10.45 4.15 10.95 8.60 ;
        RECT  10.25 7.90 10.95 8.60 ;
        RECT  11.90 3.30 12.60 4.00 ;
        RECT  12.10 3.30 12.60 10.15 ;
        RECT  12.10 9.65 14.00 10.15 ;
        RECT  13.30 9.65 14.00 10.35 ;
        RECT  13.80 4.45 14.50 5.15 ;
        RECT  14.60 5.70 15.30 6.40 ;
        RECT  12.10 5.90 15.30 6.40 ;
        RECT  15.60 3.25 16.30 3.95 ;
        RECT  13.80 4.45 16.80 4.95 ;
        RECT  15.60 7.40 16.30 8.15 ;
        RECT  15.80 3.25 16.30 9.65 ;
        RECT  15.80 8.95 16.65 9.65 ;
        RECT  15.80 4.45 16.80 5.15 ;
    END
END DFFX4
MACRO DFRRSX1
    CLASS CORE ;
    FOREIGN DFRRSX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 28.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  13.45 5.75 14.15 6.45 ;
        RECT  15.65 5.35 16.55 6.35 ;
        RECT  13.45 5.85 16.55 6.35 ;
        RECT  15.65 5.50 17.75 6.20 ;
        RECT  13.45 5.85 17.75 6.20 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  9.50 2.55 10.95 3.25 ;
        RECT  10.05 2.55 10.95 3.75 ;
        RECT  9.50 2.55 22.50 3.05 ;
        RECT  21.80 2.55 22.50 3.25 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  26.85 2.65 27.55 3.35 ;
        RECT  27.05 2.65 27.55 9.75 ;
        RECT  26.85 7.95 27.55 9.75 ;
        RECT  26.75 7.95 27.75 8.95 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  24.15 2.65 24.85 4.30 ;
        RECT  24.15 7.25 24.85 9.75 ;
        RECT  24.15 3.80 25.95 4.30 ;
        RECT  25.45 3.80 25.95 7.75 ;
        RECT  24.15 7.25 25.95 7.75 ;
        RECT  25.45 5.35 26.35 6.35 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.55 5.35 7.60 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.25 6.65 2.55 7.35 ;
        RECT  1.65 6.65 2.55 7.65 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.40 2.50 11.00 ;
        RECT  4.05 8.05 4.75 11.00 ;
        RECT  3.60 10.65 6.10 11.00 ;
        RECT  9.80 8.45 10.50 11.00 ;
        RECT  12.65 7.30 13.35 11.00 ;
        RECT  12.65 7.30 18.20 7.80 ;
        RECT  17.50 7.30 18.20 8.35 ;
        RECT  19.85 9.25 20.55 11.00 ;
        RECT  22.55 9.25 23.25 11.00 ;
        RECT  25.50 8.25 26.20 11.00 ;
        RECT  0.00 11.00 28.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.90 2.00 1.70 3.20 ;
        RECT  4.05 2.00 4.75 4.85 ;
        RECT  8.50 2.00 9.00 4.80 ;
        RECT  9.90 4.30 10.60 5.05 ;
        RECT  11.45 3.55 11.95 4.80 ;
        RECT  8.50 4.30 11.95 4.80 ;
        RECT  11.45 3.55 14.85 4.05 ;
        RECT  14.15 3.55 14.85 4.25 ;
        RECT  19.85 3.55 20.55 4.25 ;
        RECT  19.85 3.75 23.65 4.25 ;
        RECT  23.15 2.00 23.65 5.50 ;
        RECT  23.15 4.80 24.40 5.50 ;
        RECT  25.50 2.00 26.20 3.30 ;
        RECT  0.00 0.00 28.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.25 5.35 0.75 10.35 ;
        RECT  0.25 9.65 1.15 10.35 ;
        RECT  1.00 3.80 1.80 5.85 ;
        RECT  0.25 5.35 1.80 5.85 ;
        RECT  2.70 4.20 3.55 4.90 ;
        RECT  3.05 4.20 3.55 8.95 ;
        RECT  2.70 8.25 3.55 8.95 ;
        RECT  3.05 5.55 6.35 6.05 ;
        RECT  5.35 3.20 5.85 6.05 ;
        RECT  5.85 5.55 6.35 7.40 ;
        RECT  5.85 6.70 6.55 7.40 ;
        RECT  6.40 4.20 7.55 4.90 ;
        RECT  6.85 3.00 7.55 3.70 ;
        RECT  5.35 3.20 7.55 3.70 ;
        RECT  7.05 4.20 7.55 9.15 ;
        RECT  6.40 8.45 8.00 9.15 ;
        RECT  9.35 5.65 10.05 6.35 ;
        RECT  10.35 7.25 11.05 7.95 ;
        RECT  7.05 7.45 11.05 7.95 ;
        RECT  11.65 5.65 12.15 9.15 ;
        RECT  11.15 8.45 12.15 9.15 ;
        RECT  12.45 4.55 12.95 6.15 ;
        RECT  9.35 5.65 12.95 6.15 ;
        RECT  12.45 4.55 13.15 5.25 ;
        RECT  15.00 8.30 15.70 10.05 ;
        RECT  16.50 3.55 17.20 4.25 ;
        RECT  17.50 8.85 18.20 9.95 ;
        RECT  16.50 3.75 19.35 4.25 ;
        RECT  18.85 3.75 19.35 9.35 ;
        RECT  15.00 8.85 19.35 9.35 ;
        RECT  19.85 4.75 22.05 5.45 ;
        RECT  21.20 8.25 21.90 9.90 ;
        RECT  21.55 4.75 22.05 6.55 ;
        RECT  21.95 7.05 22.65 7.75 ;
        RECT  18.85 7.25 22.65 7.75 ;
        RECT  23.15 6.05 23.65 8.75 ;
        RECT  21.20 8.25 23.65 8.75 ;
        RECT  21.55 6.05 24.95 6.55 ;
        RECT  24.25 6.05 24.95 6.75 ;
    END
END DFRRSX1
MACRO DFRRSX2
    CLASS CORE ;
    FOREIGN DFRRSX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 28.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  13.45 5.75 14.15 6.45 ;
        RECT  15.65 5.35 16.55 6.35 ;
        RECT  13.45 5.85 16.55 6.35 ;
        RECT  15.65 5.50 17.75 6.20 ;
        RECT  13.45 5.85 17.75 6.20 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  9.50 2.55 10.95 3.25 ;
        RECT  10.05 2.55 10.95 3.75 ;
        RECT  9.50 2.55 22.50 3.05 ;
        RECT  21.80 2.55 22.50 3.25 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  26.85 2.65 27.55 3.35 ;
        RECT  27.05 2.65 27.55 10.50 ;
        RECT  26.85 7.95 27.55 10.50 ;
        RECT  26.75 7.95 27.75 8.95 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  24.15 2.65 24.85 4.30 ;
        RECT  24.15 7.25 24.85 10.50 ;
        RECT  24.15 3.80 25.95 4.30 ;
        RECT  25.45 3.80 25.95 7.75 ;
        RECT  24.15 7.25 25.95 7.75 ;
        RECT  25.45 5.35 26.35 6.35 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.55 5.35 7.60 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.25 6.65 2.55 7.35 ;
        RECT  1.65 6.65 2.55 7.65 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.40 2.50 11.00 ;
        RECT  4.05 8.05 4.75 11.00 ;
        RECT  3.60 10.65 6.10 11.00 ;
        RECT  9.80 8.45 10.50 11.00 ;
        RECT  12.65 7.30 13.35 11.00 ;
        RECT  12.65 7.30 18.20 7.80 ;
        RECT  17.50 7.30 18.20 8.35 ;
        RECT  19.85 9.25 20.55 11.00 ;
        RECT  22.55 9.25 23.25 11.00 ;
        RECT  25.50 8.25 26.20 11.00 ;
        RECT  0.00 11.00 28.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.90 2.00 1.70 3.20 ;
        RECT  4.05 2.00 4.75 4.85 ;
        RECT  8.50 2.00 9.00 4.80 ;
        RECT  9.90 4.30 10.60 5.05 ;
        RECT  11.45 3.55 11.95 4.80 ;
        RECT  8.50 4.30 11.95 4.80 ;
        RECT  11.45 3.55 14.85 4.05 ;
        RECT  14.15 3.55 14.85 4.25 ;
        RECT  19.85 3.55 20.55 4.25 ;
        RECT  19.85 3.75 23.65 4.25 ;
        RECT  23.15 2.00 23.65 5.50 ;
        RECT  23.15 4.80 24.40 5.50 ;
        RECT  25.50 2.00 26.20 3.30 ;
        RECT  0.00 0.00 28.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.25 5.35 0.75 10.35 ;
        RECT  0.25 9.65 1.15 10.35 ;
        RECT  1.00 3.80 1.80 5.85 ;
        RECT  0.25 5.35 1.80 5.85 ;
        RECT  2.70 4.20 3.55 4.90 ;
        RECT  3.05 4.20 3.55 8.95 ;
        RECT  2.70 8.25 3.55 8.95 ;
        RECT  3.05 5.55 6.35 6.05 ;
        RECT  5.35 3.20 5.85 6.05 ;
        RECT  5.85 5.55 6.35 7.40 ;
        RECT  5.85 6.70 6.55 7.40 ;
        RECT  6.40 4.20 7.55 4.90 ;
        RECT  6.85 3.00 7.55 3.70 ;
        RECT  5.35 3.20 7.55 3.70 ;
        RECT  7.05 4.20 7.55 9.15 ;
        RECT  6.40 8.45 8.00 9.15 ;
        RECT  9.35 5.65 10.05 6.35 ;
        RECT  10.35 7.25 11.05 7.95 ;
        RECT  7.05 7.45 11.05 7.95 ;
        RECT  11.65 5.65 12.15 9.15 ;
        RECT  11.15 8.45 12.15 9.15 ;
        RECT  12.45 4.55 12.95 6.15 ;
        RECT  9.35 5.65 12.95 6.15 ;
        RECT  12.45 4.55 13.15 5.25 ;
        RECT  15.00 8.30 15.70 10.05 ;
        RECT  16.50 3.55 17.20 4.25 ;
        RECT  17.50 8.85 18.20 9.95 ;
        RECT  16.50 3.75 19.35 4.25 ;
        RECT  18.85 3.75 19.35 9.35 ;
        RECT  15.00 8.85 19.35 9.35 ;
        RECT  19.85 4.75 22.05 5.45 ;
        RECT  21.20 8.25 21.90 9.90 ;
        RECT  21.55 4.75 22.05 6.55 ;
        RECT  21.95 7.05 22.65 7.75 ;
        RECT  18.85 7.25 22.65 7.75 ;
        RECT  23.15 6.05 23.65 8.75 ;
        RECT  21.20 8.25 23.65 8.75 ;
        RECT  21.55 6.05 24.95 6.55 ;
        RECT  24.25 6.05 24.95 6.75 ;
    END
END DFRRSX2
MACRO DFRRSX4
    CLASS CORE ;
    FOREIGN DFRRSX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 30.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  13.45 5.75 14.15 6.45 ;
        RECT  15.65 5.35 16.55 6.35 ;
        RECT  13.45 5.85 16.55 6.35 ;
        RECT  15.65 5.50 17.75 6.20 ;
        RECT  13.45 5.85 17.75 6.20 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  9.50 2.55 10.95 3.25 ;
        RECT  10.05 2.55 10.95 3.75 ;
        RECT  9.50 2.55 22.50 3.05 ;
        RECT  21.80 2.55 22.50 3.25 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  28.30 2.50 29.00 4.10 ;
        RECT  28.50 2.50 29.00 10.50 ;
        RECT  28.30 5.35 29.00 10.50 ;
        RECT  28.15 5.35 29.15 6.35 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  25.60 2.50 26.10 10.50 ;
        RECT  25.60 2.50 26.30 4.10 ;
        RECT  25.60 8.10 26.30 10.50 ;
        RECT  25.45 5.35 26.35 6.35 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.55 5.35 7.60 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.25 6.65 2.55 7.35 ;
        RECT  1.65 6.65 2.55 7.65 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.40 2.50 11.00 ;
        RECT  4.05 8.05 4.75 11.00 ;
        RECT  3.60 10.65 6.10 11.00 ;
        RECT  9.80 8.45 10.50 11.00 ;
        RECT  12.65 7.30 13.35 11.00 ;
        RECT  12.65 7.30 18.20 7.80 ;
        RECT  17.50 7.30 18.20 8.35 ;
        RECT  19.85 9.25 20.55 11.00 ;
        RECT  22.55 9.25 23.25 11.00 ;
        RECT  24.25 8.10 24.95 11.00 ;
        RECT  26.95 8.10 27.65 11.00 ;
        RECT  29.65 8.10 30.35 11.00 ;
        RECT  0.00 11.00 30.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.90 2.00 1.70 3.20 ;
        RECT  4.05 2.00 4.75 4.85 ;
        RECT  8.50 2.00 9.00 4.80 ;
        RECT  9.90 4.30 10.60 5.05 ;
        RECT  11.45 3.55 11.95 4.80 ;
        RECT  8.50 4.30 11.95 4.80 ;
        RECT  11.45 3.55 14.85 4.05 ;
        RECT  14.15 3.55 14.85 4.25 ;
        RECT  19.85 3.55 20.55 4.25 ;
        RECT  19.85 3.75 23.65 4.25 ;
        RECT  23.15 2.00 23.65 5.50 ;
        RECT  23.15 4.80 24.40 5.50 ;
        RECT  24.10 2.00 24.80 3.90 ;
        RECT  26.95 2.00 27.65 4.10 ;
        RECT  29.65 2.00 30.35 4.10 ;
        RECT  0.00 0.00 30.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.25 5.35 0.75 10.35 ;
        RECT  0.25 9.65 1.15 10.35 ;
        RECT  1.00 3.80 1.80 5.85 ;
        RECT  0.25 5.35 1.80 5.85 ;
        RECT  2.70 4.20 3.55 4.90 ;
        RECT  3.05 4.20 3.55 8.95 ;
        RECT  2.70 8.25 3.55 8.95 ;
        RECT  3.05 5.55 6.35 6.05 ;
        RECT  5.35 3.20 5.85 6.05 ;
        RECT  5.85 5.55 6.35 7.40 ;
        RECT  5.85 6.70 6.55 7.40 ;
        RECT  6.40 4.20 7.55 4.90 ;
        RECT  6.85 3.00 7.55 3.70 ;
        RECT  5.35 3.20 7.55 3.70 ;
        RECT  7.05 4.20 7.55 9.15 ;
        RECT  6.40 8.45 8.00 9.15 ;
        RECT  9.35 5.65 10.05 6.35 ;
        RECT  10.35 7.25 11.05 7.95 ;
        RECT  7.05 7.45 11.05 7.95 ;
        RECT  11.65 5.65 12.15 9.15 ;
        RECT  11.15 8.45 12.15 9.15 ;
        RECT  12.45 4.55 12.95 6.15 ;
        RECT  9.35 5.65 12.95 6.15 ;
        RECT  12.45 4.55 13.15 5.25 ;
        RECT  15.00 8.30 15.70 10.05 ;
        RECT  16.50 3.55 17.20 4.25 ;
        RECT  17.50 8.85 18.20 9.95 ;
        RECT  16.50 3.75 19.35 4.25 ;
        RECT  18.85 3.75 19.35 9.35 ;
        RECT  15.00 8.85 19.35 9.35 ;
        RECT  19.85 4.75 22.05 5.45 ;
        RECT  21.20 8.25 21.90 9.90 ;
        RECT  21.55 4.75 22.05 6.55 ;
        RECT  21.95 7.05 22.65 7.75 ;
        RECT  18.85 7.25 22.65 7.75 ;
        RECT  23.15 6.05 23.65 8.75 ;
        RECT  21.20 8.25 23.65 8.75 ;
        RECT  21.55 6.05 24.95 6.55 ;
        RECT  24.25 6.05 24.95 6.75 ;
    END
END DFRRSX4
MACRO DFRRX1
    CLASS CORE ;
    FOREIGN DFRRX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 25.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  9.50 2.55 10.20 3.25 ;
        RECT  15.65 2.55 16.55 3.75 ;
        RECT  9.50 2.55 19.70 3.05 ;
        RECT  19.00 2.55 19.70 3.25 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  24.05 2.65 24.75 3.35 ;
        RECT  24.25 2.65 24.75 9.75 ;
        RECT  24.05 7.95 24.75 9.75 ;
        RECT  23.95 7.95 24.95 8.95 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  21.35 2.65 22.05 4.30 ;
        RECT  21.35 7.25 22.05 9.75 ;
        RECT  21.35 3.80 23.15 4.30 ;
        RECT  22.65 3.80 23.15 7.75 ;
        RECT  21.35 7.25 23.15 7.75 ;
        RECT  22.65 5.35 23.55 6.35 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.55 5.35 7.60 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.25 6.65 2.55 7.35 ;
        RECT  1.65 6.65 2.55 7.65 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.40 2.50 11.00 ;
        RECT  4.05 8.05 4.75 11.00 ;
        RECT  9.80 8.20 10.50 11.00 ;
        RECT  12.30 9.55 13.00 11.00 ;
        RECT  17.15 9.30 17.85 11.00 ;
        RECT  19.85 9.30 20.55 11.00 ;
        RECT  22.70 8.25 23.40 11.00 ;
        RECT  0.00 11.00 25.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.90 2.00 1.70 3.20 ;
        RECT  4.05 2.00 4.75 4.85 ;
        RECT  8.50 2.00 9.00 4.25 ;
        RECT  9.90 3.75 10.60 4.95 ;
        RECT  8.50 3.75 13.60 4.25 ;
        RECT  12.90 3.75 13.60 5.45 ;
        RECT  18.55 3.75 19.25 5.45 ;
        RECT  17.60 4.70 19.25 5.45 ;
        RECT  20.35 2.00 20.85 4.25 ;
        RECT  18.55 3.75 20.85 4.25 ;
        RECT  22.70 2.00 23.40 3.30 ;
        RECT  0.00 0.00 25.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  16.95 6.05 22.15 6.50 ;
        RECT  0.25 5.35 0.75 10.35 ;
        RECT  0.25 9.65 1.15 10.35 ;
        RECT  1.00 3.80 1.80 5.85 ;
        RECT  0.25 5.35 1.80 5.85 ;
        RECT  2.70 4.20 3.55 4.90 ;
        RECT  3.05 4.20 3.55 8.95 ;
        RECT  2.70 8.25 3.55 8.95 ;
        RECT  3.05 5.55 6.35 6.05 ;
        RECT  5.35 3.20 5.85 6.05 ;
        RECT  5.85 5.55 6.35 7.40 ;
        RECT  5.85 6.70 6.55 7.40 ;
        RECT  6.40 4.20 7.55 4.90 ;
        RECT  6.85 3.00 7.55 3.70 ;
        RECT  5.35 3.20 7.55 3.70 ;
        RECT  7.05 4.20 7.55 9.25 ;
        RECT  6.40 8.55 8.00 9.25 ;
        RECT  9.35 5.65 10.05 6.35 ;
        RECT  10.35 6.90 11.05 7.60 ;
        RECT  7.05 7.10 11.05 7.60 ;
        RECT  11.40 4.75 12.10 6.15 ;
        RECT  9.35 5.65 12.10 6.15 ;
        RECT  11.60 4.75 12.10 8.85 ;
        RECT  11.15 8.10 12.10 8.85 ;
        RECT  15.25 4.75 15.50 10.05 ;
        RECT  14.80 7.30 15.50 10.05 ;
        RECT  15.25 4.75 15.75 7.80 ;
        RECT  15.25 4.75 15.95 5.45 ;
        RECT  16.95 6.00 17.65 6.70 ;
        RECT  18.50 8.30 19.20 9.95 ;
        RECT  19.15 7.10 19.85 7.80 ;
        RECT  14.80 7.30 19.85 7.80 ;
        RECT  20.35 6.00 20.85 8.80 ;
        RECT  18.50 8.30 20.85 8.80 ;
        RECT  20.90 4.80 21.60 6.75 ;
        RECT  16.95 6.00 21.60 6.50 ;
        RECT  20.35 6.05 22.15 6.75 ;
    END
END DFRRX1
MACRO DFRRX2
    CLASS CORE ;
    FOREIGN DFRRX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 25.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  9.50 2.55 10.20 3.25 ;
        RECT  15.65 2.55 16.55 3.75 ;
        RECT  9.50 2.55 19.70 3.05 ;
        RECT  19.00 2.55 19.70 3.25 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  24.05 2.65 24.75 3.35 ;
        RECT  24.25 2.65 24.75 10.50 ;
        RECT  24.05 7.95 24.75 10.50 ;
        RECT  23.95 7.95 24.95 8.95 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  21.35 2.65 22.05 4.30 ;
        RECT  21.35 7.25 22.05 10.50 ;
        RECT  21.35 3.80 23.15 4.30 ;
        RECT  22.65 3.80 23.15 7.75 ;
        RECT  21.35 7.25 23.15 7.75 ;
        RECT  22.65 5.35 23.55 6.35 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.55 5.35 7.60 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.25 6.65 2.55 7.35 ;
        RECT  1.65 6.65 2.55 7.65 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.40 2.50 11.00 ;
        RECT  4.05 8.05 4.75 11.00 ;
        RECT  9.80 8.20 10.50 11.00 ;
        RECT  12.30 9.55 13.00 11.00 ;
        RECT  17.15 9.30 17.85 11.00 ;
        RECT  19.85 9.30 20.55 11.00 ;
        RECT  22.70 8.25 23.40 11.00 ;
        RECT  0.00 11.00 25.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.90 2.00 1.70 3.20 ;
        RECT  4.05 2.00 4.75 4.85 ;
        RECT  8.50 2.00 9.00 4.25 ;
        RECT  9.90 3.75 10.60 4.95 ;
        RECT  8.50 3.75 13.60 4.25 ;
        RECT  12.90 3.75 13.60 5.45 ;
        RECT  18.55 3.75 19.25 5.45 ;
        RECT  17.60 4.70 19.25 5.45 ;
        RECT  20.35 2.00 20.85 4.25 ;
        RECT  18.55 3.75 20.85 4.25 ;
        RECT  22.70 2.00 23.40 3.30 ;
        RECT  0.00 0.00 25.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  16.95 6.05 22.15 6.50 ;
        RECT  0.25 5.35 0.75 10.35 ;
        RECT  0.25 9.65 1.15 10.35 ;
        RECT  1.00 3.80 1.80 5.85 ;
        RECT  0.25 5.35 1.80 5.85 ;
        RECT  2.70 4.20 3.55 4.90 ;
        RECT  3.05 4.20 3.55 8.95 ;
        RECT  2.70 8.25 3.55 8.95 ;
        RECT  3.05 5.55 6.35 6.05 ;
        RECT  5.35 3.20 5.85 6.05 ;
        RECT  5.85 5.55 6.35 7.40 ;
        RECT  5.85 6.70 6.55 7.40 ;
        RECT  6.40 4.20 7.55 4.90 ;
        RECT  6.85 3.00 7.55 3.70 ;
        RECT  5.35 3.20 7.55 3.70 ;
        RECT  7.05 4.20 7.55 9.25 ;
        RECT  6.40 8.55 8.00 9.25 ;
        RECT  9.35 5.65 10.05 6.35 ;
        RECT  10.35 6.90 11.05 7.60 ;
        RECT  7.05 7.10 11.05 7.60 ;
        RECT  11.40 4.75 12.10 6.15 ;
        RECT  9.35 5.65 12.10 6.15 ;
        RECT  11.60 4.75 12.10 8.85 ;
        RECT  11.15 8.10 12.10 8.85 ;
        RECT  15.25 4.75 15.50 10.05 ;
        RECT  14.80 7.30 15.50 10.05 ;
        RECT  15.25 4.75 15.75 7.80 ;
        RECT  15.25 4.75 15.95 5.45 ;
        RECT  16.95 6.00 17.65 6.70 ;
        RECT  18.50 8.30 19.20 9.95 ;
        RECT  19.15 7.10 19.85 7.80 ;
        RECT  14.80 7.30 19.85 7.80 ;
        RECT  20.35 6.00 20.85 8.80 ;
        RECT  18.50 8.30 20.85 8.80 ;
        RECT  20.90 4.80 21.60 6.75 ;
        RECT  16.95 6.00 21.60 6.50 ;
        RECT  20.35 6.05 22.15 6.75 ;
    END
END DFRRX2
MACRO DFRRX4
    CLASS CORE ;
    FOREIGN DFRRX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 28.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  9.50 2.55 10.20 3.25 ;
        RECT  15.65 2.55 16.55 3.75 ;
        RECT  9.50 2.55 19.70 3.05 ;
        RECT  19.00 2.55 19.70 3.25 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  25.50 2.50 26.20 4.10 ;
        RECT  25.70 2.50 26.20 10.50 ;
        RECT  25.50 5.35 26.20 10.50 ;
        RECT  25.35 5.35 26.35 6.35 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  22.80 2.50 23.30 10.50 ;
        RECT  22.80 2.50 23.50 4.10 ;
        RECT  22.80 8.10 23.50 10.50 ;
        RECT  22.65 5.35 23.55 6.35 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.55 5.35 7.60 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.25 6.65 2.55 7.35 ;
        RECT  1.65 6.65 2.55 7.65 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.40 2.50 11.00 ;
        RECT  4.05 8.05 4.75 11.00 ;
        RECT  9.80 8.20 10.50 11.00 ;
        RECT  12.30 9.55 13.00 11.00 ;
        RECT  17.15 9.30 17.85 11.00 ;
        RECT  19.85 9.30 20.55 11.00 ;
        RECT  21.45 8.10 22.15 11.00 ;
        RECT  24.15 8.10 24.85 11.00 ;
        RECT  26.85 8.10 27.55 11.00 ;
        RECT  0.00 11.00 28.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.90 2.00 1.70 3.20 ;
        RECT  4.05 2.00 4.75 4.85 ;
        RECT  8.50 2.00 9.00 4.25 ;
        RECT  9.90 3.75 10.60 4.95 ;
        RECT  8.50 3.75 13.60 4.25 ;
        RECT  12.90 3.75 13.60 5.45 ;
        RECT  18.55 3.75 19.25 5.45 ;
        RECT  17.60 4.70 19.25 5.45 ;
        RECT  21.30 2.00 22.00 4.25 ;
        RECT  18.55 3.75 22.00 4.25 ;
        RECT  24.15 2.00 24.85 4.10 ;
        RECT  26.85 2.00 27.55 4.10 ;
        RECT  0.00 0.00 28.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.25 5.35 0.75 10.35 ;
        RECT  0.25 9.65 1.15 10.35 ;
        RECT  1.00 3.80 1.80 5.85 ;
        RECT  0.25 5.35 1.80 5.85 ;
        RECT  2.70 4.20 3.55 4.90 ;
        RECT  3.05 4.20 3.55 8.95 ;
        RECT  2.70 8.25 3.55 8.95 ;
        RECT  3.05 5.55 6.35 6.05 ;
        RECT  5.35 3.20 5.85 6.05 ;
        RECT  5.85 5.55 6.35 7.40 ;
        RECT  5.85 6.70 6.55 7.40 ;
        RECT  6.40 4.20 7.55 4.90 ;
        RECT  6.85 3.00 7.55 3.70 ;
        RECT  5.35 3.20 7.55 3.70 ;
        RECT  7.05 4.20 7.55 9.25 ;
        RECT  6.40 8.55 8.00 9.25 ;
        RECT  9.35 5.65 10.05 6.35 ;
        RECT  10.35 6.90 11.05 7.60 ;
        RECT  7.05 7.10 11.05 7.60 ;
        RECT  11.40 4.75 12.10 6.15 ;
        RECT  9.35 5.65 12.10 6.15 ;
        RECT  11.60 4.75 12.10 8.85 ;
        RECT  11.15 8.10 12.10 8.85 ;
        RECT  15.25 4.75 15.50 10.05 ;
        RECT  14.80 7.30 15.50 10.05 ;
        RECT  15.25 4.75 15.75 7.80 ;
        RECT  15.25 4.75 15.95 5.45 ;
        RECT  16.95 6.00 17.65 6.70 ;
        RECT  18.50 8.30 19.20 9.95 ;
        RECT  19.15 7.10 19.85 7.80 ;
        RECT  14.80 7.30 19.85 7.80 ;
        RECT  20.35 6.00 20.85 8.80 ;
        RECT  18.50 8.30 20.85 8.80 ;
        RECT  16.95 6.00 22.15 6.50 ;
        RECT  21.45 4.75 21.65 6.70 ;
        RECT  20.95 4.75 21.65 6.50 ;
        RECT  21.45 6.00 22.15 6.70 ;
    END
END DFRRX4
MACRO DFRSX1
    CLASS CORE ;
    FOREIGN DFRSX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  11.45 7.05 12.15 8.40 ;
        RECT  12.85 6.70 13.75 7.60 ;
        RECT  13.25 5.45 13.75 7.60 ;
        RECT  11.45 7.05 13.75 7.60 ;
        RECT  13.90 5.25 14.60 5.95 ;
        RECT  13.25 5.45 14.60 5.95 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  19.95 3.75 20.65 4.45 ;
        RECT  20.10 3.75 20.65 8.85 ;
        RECT  19.95 7.15 20.65 8.85 ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  22.65 3.75 23.35 4.45 ;
        RECT  22.85 3.75 23.35 8.85 ;
        RECT  22.65 7.15 23.35 8.85 ;
        RECT  22.65 5.40 23.55 6.30 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.55 5.35 7.60 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.25 6.65 2.55 7.35 ;
        RECT  1.65 6.65 2.55 7.65 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.40 2.50 11.00 ;
        RECT  4.05 8.05 4.75 11.00 ;
        RECT  3.40 10.65 6.95 11.00 ;
        RECT  8.75 7.90 9.45 11.00 ;
        RECT  8.00 10.60 9.60 11.00 ;
        RECT  12.05 8.90 12.75 11.00 ;
        RECT  17.05 7.40 17.75 11.00 ;
        RECT  21.30 7.15 22.00 11.00 ;
        RECT  17.05 10.70 23.35 11.00 ;
        RECT  0.00 11.00 23.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.90 2.00 1.70 3.20 ;
        RECT  4.05 2.00 4.75 4.85 ;
        RECT  8.15 2.00 9.75 3.15 ;
        RECT  9.05 2.00 9.75 4.90 ;
        RECT  11.20 2.00 11.90 3.25 ;
        RECT  17.05 2.00 17.75 3.95 ;
        RECT  21.30 2.00 22.00 4.45 ;
        RECT  0.00 0.00 23.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.25 5.35 0.75 10.35 ;
        RECT  0.25 9.65 1.20 10.35 ;
        RECT  1.00 3.80 1.80 5.85 ;
        RECT  0.25 5.35 1.80 5.85 ;
        RECT  2.70 4.20 3.55 4.90 ;
        RECT  3.05 4.20 3.55 8.95 ;
        RECT  2.70 8.25 3.55 8.95 ;
        RECT  3.05 5.55 6.35 6.05 ;
        RECT  5.35 3.20 5.85 6.05 ;
        RECT  5.85 5.55 6.35 7.40 ;
        RECT  5.85 6.70 6.55 7.40 ;
        RECT  6.40 4.20 7.10 4.90 ;
        RECT  6.40 4.40 7.55 4.90 ;
        RECT  7.05 4.20 7.10 9.55 ;
        RECT  6.40 7.90 7.10 9.55 ;
        RECT  6.85 3.00 7.55 3.70 ;
        RECT  5.35 3.20 7.55 3.70 ;
        RECT  7.05 4.40 7.55 8.40 ;
        RECT  6.40 7.90 7.55 8.40 ;
        RECT  8.30 5.45 9.00 6.15 ;
        RECT  7.05 6.70 9.95 7.20 ;
        RECT  9.25 6.70 9.95 7.40 ;
        RECT  8.30 5.45 10.95 5.95 ;
        RECT  10.45 4.35 10.95 9.55 ;
        RECT  10.45 8.85 11.25 9.55 ;
        RECT  11.55 4.15 12.25 4.85 ;
        RECT  10.45 4.35 12.25 4.85 ;
        RECT  13.70 3.30 14.40 4.00 ;
        RECT  13.70 3.45 15.60 4.00 ;
        RECT  14.55 7.20 15.10 10.50 ;
        RECT  14.40 8.75 15.10 10.50 ;
        RECT  15.10 3.45 15.60 7.90 ;
        RECT  14.55 7.20 15.60 7.90 ;
        RECT  16.60 4.45 17.30 5.15 ;
        RECT  17.40 5.70 18.10 6.40 ;
        RECT  15.10 5.90 18.10 6.40 ;
        RECT  18.40 3.25 19.10 3.95 ;
        RECT  16.60 4.45 19.10 4.95 ;
        RECT  18.60 3.25 19.10 10.10 ;
        RECT  18.40 7.40 19.10 10.10 ;
    END
END DFRSX1
MACRO DFRSX2
    CLASS CORE ;
    FOREIGN DFRSX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  11.45 7.05 12.15 8.40 ;
        RECT  12.85 6.70 13.75 7.60 ;
        RECT  13.25 5.45 13.75 7.60 ;
        RECT  11.45 7.05 13.75 7.60 ;
        RECT  13.90 5.25 14.60 5.95 ;
        RECT  13.25 5.45 14.60 5.95 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  19.95 2.70 20.65 4.50 ;
        RECT  20.10 2.70 20.65 10.50 ;
        RECT  19.95 7.10 20.65 10.50 ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  22.65 2.70 23.35 4.50 ;
        RECT  22.85 2.70 23.35 10.50 ;
        RECT  22.65 7.10 23.35 10.50 ;
        RECT  22.65 5.40 23.55 6.30 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.55 5.35 7.60 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.25 6.65 2.55 7.35 ;
        RECT  1.65 6.65 2.55 7.65 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.40 2.50 11.00 ;
        RECT  4.05 8.05 4.75 11.00 ;
        RECT  3.40 10.65 6.95 11.00 ;
        RECT  8.75 7.90 9.45 11.00 ;
        RECT  8.00 10.60 9.60 11.00 ;
        RECT  12.05 8.90 12.75 11.00 ;
        RECT  17.05 7.40 17.75 11.00 ;
        RECT  21.30 7.10 22.00 11.00 ;
        RECT  0.00 11.00 23.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.90 2.00 1.70 3.20 ;
        RECT  4.05 2.00 4.75 4.85 ;
        RECT  8.15 2.00 9.75 3.15 ;
        RECT  9.05 2.00 9.75 4.90 ;
        RECT  11.20 2.00 11.90 3.25 ;
        RECT  17.05 2.00 17.75 3.95 ;
        RECT  21.30 2.00 22.00 4.50 ;
        RECT  0.00 0.00 23.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.25 5.35 0.75 10.35 ;
        RECT  0.25 9.65 1.20 10.35 ;
        RECT  1.00 3.80 1.80 5.85 ;
        RECT  0.25 5.35 1.80 5.85 ;
        RECT  2.70 4.20 3.55 4.90 ;
        RECT  3.05 4.20 3.55 8.95 ;
        RECT  2.70 8.25 3.55 8.95 ;
        RECT  3.05 5.55 6.35 6.05 ;
        RECT  5.35 3.20 5.85 6.05 ;
        RECT  5.85 5.55 6.35 7.40 ;
        RECT  5.85 6.70 6.55 7.40 ;
        RECT  6.40 4.20 7.10 4.90 ;
        RECT  6.40 4.40 7.55 4.90 ;
        RECT  7.05 4.20 7.10 9.55 ;
        RECT  6.40 7.90 7.10 9.55 ;
        RECT  6.85 3.00 7.55 3.70 ;
        RECT  5.35 3.20 7.55 3.70 ;
        RECT  7.05 4.40 7.55 8.40 ;
        RECT  6.40 7.90 7.55 8.40 ;
        RECT  8.30 5.45 9.00 6.15 ;
        RECT  7.05 6.70 9.95 7.20 ;
        RECT  9.25 6.70 9.95 7.40 ;
        RECT  8.30 5.45 10.95 5.95 ;
        RECT  10.45 4.35 10.95 9.55 ;
        RECT  10.45 8.85 11.25 9.55 ;
        RECT  11.55 4.15 12.25 4.85 ;
        RECT  10.45 4.35 12.25 4.85 ;
        RECT  13.70 3.30 14.40 4.00 ;
        RECT  13.70 3.45 15.60 4.00 ;
        RECT  14.55 7.20 15.10 10.50 ;
        RECT  14.40 8.75 15.10 10.50 ;
        RECT  15.10 3.45 15.60 7.90 ;
        RECT  14.55 7.20 15.60 7.90 ;
        RECT  16.60 4.45 17.30 5.15 ;
        RECT  17.40 5.70 18.10 6.40 ;
        RECT  15.10 5.90 18.10 6.40 ;
        RECT  18.40 3.25 19.10 3.95 ;
        RECT  16.60 4.45 19.10 4.95 ;
        RECT  18.60 3.25 19.10 10.10 ;
        RECT  18.40 7.40 19.10 10.10 ;
    END
END DFRSX2
MACRO DFRSX4
    CLASS CORE ;
    FOREIGN DFRSX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 26.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  11.45 7.05 12.15 8.40 ;
        RECT  12.85 6.70 13.75 7.60 ;
        RECT  13.25 5.45 13.75 7.60 ;
        RECT  11.45 7.05 13.75 7.60 ;
        RECT  13.90 5.25 14.60 5.95 ;
        RECT  13.25 5.45 14.60 5.95 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  21.40 2.70 21.90 10.50 ;
        RECT  21.40 2.70 22.10 4.50 ;
        RECT  21.40 7.10 22.10 10.50 ;
        RECT  21.25 5.35 22.15 6.35 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  24.10 2.70 24.80 4.50 ;
        RECT  24.30 2.70 24.80 10.50 ;
        RECT  24.10 5.35 24.80 10.50 ;
        RECT  23.95 5.35 24.95 6.35 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.55 5.35 7.60 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.25 6.65 2.55 7.35 ;
        RECT  1.65 6.65 2.55 7.65 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.40 2.50 11.00 ;
        RECT  4.05 8.05 4.75 11.00 ;
        RECT  3.40 10.65 6.95 11.00 ;
        RECT  8.75 7.90 9.45 11.00 ;
        RECT  8.00 10.60 9.60 11.00 ;
        RECT  12.05 8.90 12.75 11.00 ;
        RECT  17.05 7.40 17.75 11.00 ;
        RECT  20.05 7.10 20.75 11.00 ;
        RECT  22.75 7.10 23.45 11.00 ;
        RECT  25.45 7.10 26.15 11.00 ;
        RECT  0.00 11.00 26.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.90 2.00 1.70 3.20 ;
        RECT  4.05 2.00 4.75 4.85 ;
        RECT  8.15 2.00 9.75 3.15 ;
        RECT  9.05 2.00 9.75 4.90 ;
        RECT  11.20 2.00 11.90 3.25 ;
        RECT  17.05 2.00 17.75 3.95 ;
        RECT  20.05 2.00 20.75 4.50 ;
        RECT  22.75 2.00 23.45 4.50 ;
        RECT  25.45 2.00 26.15 4.50 ;
        RECT  0.00 0.00 26.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.25 5.35 0.75 10.35 ;
        RECT  0.25 9.65 1.20 10.35 ;
        RECT  1.00 3.80 1.80 5.85 ;
        RECT  0.25 5.35 1.80 5.85 ;
        RECT  2.70 4.20 3.55 4.90 ;
        RECT  3.05 4.20 3.55 8.95 ;
        RECT  2.70 8.25 3.55 8.95 ;
        RECT  3.05 5.55 6.35 6.05 ;
        RECT  5.35 3.20 5.85 6.05 ;
        RECT  5.85 5.55 6.35 7.40 ;
        RECT  5.85 6.70 6.55 7.40 ;
        RECT  6.40 4.20 7.10 4.90 ;
        RECT  6.40 4.40 7.55 4.90 ;
        RECT  7.05 4.20 7.10 9.55 ;
        RECT  6.40 7.90 7.10 9.55 ;
        RECT  6.85 3.00 7.55 3.70 ;
        RECT  5.35 3.20 7.55 3.70 ;
        RECT  7.05 4.40 7.55 8.40 ;
        RECT  6.40 7.90 7.55 8.40 ;
        RECT  8.30 5.45 9.00 6.15 ;
        RECT  7.05 6.70 9.95 7.20 ;
        RECT  9.25 6.70 9.95 7.40 ;
        RECT  8.30 5.45 10.95 5.95 ;
        RECT  10.45 4.35 10.95 9.55 ;
        RECT  10.45 8.85 11.25 9.55 ;
        RECT  11.55 4.15 12.25 4.85 ;
        RECT  10.45 4.35 12.25 4.85 ;
        RECT  13.70 3.30 14.40 4.00 ;
        RECT  13.70 3.45 15.60 4.00 ;
        RECT  14.55 7.20 15.10 10.50 ;
        RECT  14.40 8.75 15.10 10.50 ;
        RECT  15.10 3.45 15.60 7.90 ;
        RECT  14.55 7.20 15.60 7.90 ;
        RECT  16.60 4.45 17.30 5.15 ;
        RECT  17.40 5.70 18.10 6.40 ;
        RECT  15.10 5.90 18.10 6.40 ;
        RECT  18.40 3.25 19.10 3.95 ;
        RECT  16.60 4.45 19.10 4.95 ;
        RECT  18.60 3.25 19.10 10.10 ;
        RECT  18.40 7.40 19.10 10.10 ;
    END
END DFRSX4
MACRO DFRX1
    CLASS CORE ;
    FOREIGN DFRX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  17.15 3.75 17.85 4.45 ;
        RECT  17.30 3.75 17.85 8.85 ;
        RECT  17.15 7.15 17.85 8.85 ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  19.85 3.75 20.55 4.45 ;
        RECT  20.05 3.75 20.55 8.85 ;
        RECT  19.85 7.15 20.55 8.85 ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.55 5.35 7.60 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.25 6.65 2.55 7.35 ;
        RECT  1.65 6.65 2.55 7.65 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.40 2.50 11.00 ;
        RECT  4.05 8.05 4.75 11.00 ;
        RECT  3.40 10.65 6.95 11.00 ;
        RECT  8.75 7.90 9.45 11.00 ;
        RECT  8.00 10.45 10.15 11.00 ;
        RECT  10.95 10.40 11.65 11.00 ;
        RECT  14.25 7.40 14.95 8.15 ;
        RECT  14.45 7.40 14.95 11.00 ;
        RECT  15.80 10.15 16.50 11.00 ;
        RECT  18.50 7.15 19.20 11.00 ;
        RECT  17.30 10.70 20.55 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.90 2.00 1.70 3.20 ;
        RECT  4.05 2.00 4.75 4.85 ;
        RECT  8.75 2.00 9.45 4.90 ;
        RECT  8.75 2.00 10.10 3.10 ;
        RECT  14.25 2.00 14.95 3.95 ;
        RECT  18.50 2.00 19.20 4.45 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.25 5.35 0.75 10.35 ;
        RECT  0.25 9.65 1.20 10.35 ;
        RECT  1.00 3.80 1.80 5.85 ;
        RECT  0.25 5.35 1.80 5.85 ;
        RECT  2.70 4.20 3.55 4.90 ;
        RECT  3.05 4.20 3.55 8.95 ;
        RECT  2.70 8.25 3.55 8.95 ;
        RECT  3.05 5.55 6.35 6.05 ;
        RECT  5.35 3.20 5.85 6.05 ;
        RECT  5.85 5.55 6.35 7.40 ;
        RECT  5.85 6.70 6.55 7.40 ;
        RECT  6.40 4.20 7.10 4.90 ;
        RECT  6.40 4.40 7.55 4.90 ;
        RECT  7.05 4.20 7.10 9.55 ;
        RECT  6.40 7.90 7.10 9.55 ;
        RECT  6.85 3.00 7.55 3.70 ;
        RECT  5.35 3.20 7.55 3.70 ;
        RECT  7.05 4.40 7.55 8.40 ;
        RECT  6.40 7.90 7.55 8.40 ;
        RECT  8.30 5.45 9.00 6.15 ;
        RECT  7.05 6.70 9.95 7.20 ;
        RECT  9.25 6.70 9.95 7.40 ;
        RECT  8.30 5.45 10.95 5.95 ;
        RECT  10.45 4.15 10.80 8.60 ;
        RECT  10.10 4.15 10.80 5.95 ;
        RECT  10.45 5.45 10.95 8.60 ;
        RECT  10.25 7.90 10.95 8.60 ;
        RECT  11.75 2.45 12.60 3.15 ;
        RECT  11.90 2.45 12.60 4.05 ;
        RECT  12.10 2.45 12.60 10.15 ;
        RECT  12.10 9.65 14.00 10.15 ;
        RECT  13.30 9.65 14.00 10.35 ;
        RECT  13.80 4.45 14.50 5.15 ;
        RECT  14.60 5.70 15.30 6.40 ;
        RECT  12.10 5.90 15.30 6.40 ;
        RECT  15.60 3.25 16.30 3.95 ;
        RECT  13.80 4.45 16.30 4.95 ;
        RECT  15.60 7.40 16.30 8.15 ;
        RECT  15.80 3.25 16.30 9.65 ;
        RECT  15.80 8.95 16.65 9.65 ;
    END
END DFRX1
MACRO DFRX2
    CLASS CORE ;
    FOREIGN DFRX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  17.15 2.70 17.85 4.50 ;
        RECT  17.30 2.70 17.85 9.60 ;
        RECT  17.15 7.10 17.85 9.60 ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  19.85 2.70 20.55 4.50 ;
        RECT  20.05 2.70 20.55 10.50 ;
        RECT  19.85 7.10 20.55 10.50 ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.55 5.35 7.60 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.25 6.65 2.55 7.35 ;
        RECT  1.65 6.65 2.55 7.65 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.40 2.50 11.00 ;
        RECT  4.05 8.05 4.75 11.00 ;
        RECT  3.40 10.65 6.95 11.00 ;
        RECT  8.75 7.90 9.45 11.00 ;
        RECT  8.00 10.45 10.15 11.00 ;
        RECT  10.95 10.40 11.65 11.00 ;
        RECT  14.25 7.40 14.95 8.15 ;
        RECT  14.45 7.40 14.95 11.00 ;
        RECT  15.80 10.20 16.50 11.00 ;
        RECT  18.50 7.10 19.20 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.90 2.00 1.70 3.20 ;
        RECT  4.05 2.00 4.75 4.85 ;
        RECT  8.75 2.00 9.45 4.90 ;
        RECT  8.75 2.00 10.10 3.10 ;
        RECT  14.25 2.00 14.95 4.00 ;
        RECT  18.50 2.00 19.20 4.50 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.25 5.35 0.75 10.35 ;
        RECT  0.25 9.65 1.20 10.35 ;
        RECT  1.00 3.80 1.80 5.85 ;
        RECT  0.25 5.35 1.80 5.85 ;
        RECT  2.70 4.20 3.55 4.90 ;
        RECT  3.05 4.20 3.55 8.95 ;
        RECT  2.70 8.25 3.55 8.95 ;
        RECT  3.05 5.55 6.35 6.05 ;
        RECT  5.35 3.20 5.85 6.05 ;
        RECT  5.85 5.55 6.35 7.40 ;
        RECT  5.85 6.70 6.55 7.40 ;
        RECT  6.40 4.20 7.10 4.90 ;
        RECT  6.40 4.40 7.55 4.90 ;
        RECT  7.05 4.20 7.10 9.55 ;
        RECT  6.40 7.90 7.10 9.55 ;
        RECT  6.85 3.00 7.55 3.70 ;
        RECT  5.35 3.20 7.55 3.70 ;
        RECT  7.05 4.40 7.55 8.40 ;
        RECT  6.40 7.90 7.55 8.40 ;
        RECT  8.30 5.45 9.00 6.15 ;
        RECT  7.05 6.70 9.95 7.20 ;
        RECT  9.25 6.70 9.95 7.40 ;
        RECT  8.30 5.45 10.95 5.95 ;
        RECT  10.45 4.15 10.80 8.60 ;
        RECT  10.10 4.15 10.80 5.95 ;
        RECT  10.45 5.45 10.95 8.60 ;
        RECT  10.25 7.90 10.95 8.60 ;
        RECT  11.75 2.45 12.60 3.15 ;
        RECT  11.90 2.45 12.60 4.05 ;
        RECT  12.10 2.45 12.60 10.15 ;
        RECT  12.10 9.65 14.00 10.15 ;
        RECT  13.30 9.65 14.00 10.35 ;
        RECT  13.80 4.45 14.50 5.15 ;
        RECT  14.60 5.70 15.30 6.40 ;
        RECT  12.10 5.90 15.30 6.40 ;
        RECT  15.60 3.30 16.30 4.95 ;
        RECT  13.80 4.45 16.30 4.95 ;
        RECT  15.60 7.40 16.30 8.15 ;
        RECT  15.80 3.30 16.30 9.65 ;
        RECT  15.80 8.95 16.65 9.65 ;
    END
END DFRX2
MACRO DFRX4
    CLASS CORE ;
    FOREIGN DFRX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  18.60 2.70 19.10 10.50 ;
        RECT  18.60 2.70 19.30 4.50 ;
        RECT  18.60 7.10 19.30 10.50 ;
        RECT  18.45 5.35 19.35 6.35 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  21.30 2.70 22.00 4.50 ;
        RECT  21.50 2.70 22.00 10.50 ;
        RECT  21.30 5.35 22.00 10.50 ;
        RECT  21.15 5.35 22.15 6.35 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.55 5.35 7.60 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.25 6.65 2.55 7.35 ;
        RECT  1.65 6.65 2.55 7.65 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.40 2.50 11.00 ;
        RECT  4.05 8.05 4.75 11.00 ;
        RECT  3.40 10.65 6.95 11.00 ;
        RECT  8.75 7.90 9.45 11.00 ;
        RECT  8.00 10.45 10.10 11.00 ;
        RECT  10.90 10.40 11.60 11.00 ;
        RECT  14.25 7.40 14.95 8.15 ;
        RECT  14.45 7.40 14.95 11.00 ;
        RECT  15.75 10.15 16.45 11.00 ;
        RECT  17.25 7.10 17.95 11.00 ;
        RECT  19.95 7.10 20.65 11.00 ;
        RECT  22.65 7.10 23.35 11.00 ;
        RECT  0.00 11.00 23.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.90 2.00 1.70 3.20 ;
        RECT  4.05 2.00 4.75 4.85 ;
        RECT  8.75 2.00 9.45 4.90 ;
        RECT  8.75 2.00 10.10 3.10 ;
        RECT  14.25 2.00 14.95 3.95 ;
        RECT  17.25 2.00 17.95 4.50 ;
        RECT  19.95 2.00 20.65 4.50 ;
        RECT  22.65 2.00 23.35 4.50 ;
        RECT  0.00 0.00 23.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.25 5.35 0.75 10.35 ;
        RECT  0.25 9.65 1.20 10.35 ;
        RECT  1.00 3.80 1.80 5.85 ;
        RECT  0.25 5.35 1.80 5.85 ;
        RECT  2.70 4.20 3.55 4.90 ;
        RECT  3.05 4.20 3.55 8.95 ;
        RECT  2.70 8.25 3.55 8.95 ;
        RECT  3.05 5.55 6.35 6.05 ;
        RECT  5.35 3.20 5.85 6.05 ;
        RECT  5.85 5.55 6.35 7.40 ;
        RECT  5.85 6.70 6.55 7.40 ;
        RECT  6.40 4.20 7.10 4.90 ;
        RECT  6.40 4.40 7.55 4.90 ;
        RECT  7.05 4.20 7.10 9.55 ;
        RECT  6.40 7.90 7.10 9.55 ;
        RECT  6.85 3.00 7.55 3.70 ;
        RECT  5.35 3.20 7.55 3.70 ;
        RECT  7.05 4.40 7.55 8.40 ;
        RECT  6.40 7.90 7.55 8.40 ;
        RECT  8.30 5.45 9.00 6.15 ;
        RECT  7.05 6.70 9.95 7.20 ;
        RECT  9.25 6.70 9.95 7.40 ;
        RECT  8.30 5.45 10.95 5.95 ;
        RECT  10.45 4.15 10.80 8.60 ;
        RECT  10.10 4.15 10.80 5.95 ;
        RECT  10.45 5.45 10.95 8.60 ;
        RECT  10.25 7.90 10.95 8.60 ;
        RECT  11.75 2.45 12.60 3.15 ;
        RECT  11.90 2.45 12.60 4.05 ;
        RECT  12.10 2.45 12.60 10.15 ;
        RECT  12.10 9.65 13.95 10.15 ;
        RECT  13.25 9.65 13.95 10.35 ;
        RECT  13.80 4.45 14.50 5.15 ;
        RECT  14.60 5.70 15.30 6.40 ;
        RECT  12.10 5.90 15.30 6.40 ;
        RECT  15.60 3.25 16.30 3.95 ;
        RECT  13.80 4.45 16.30 4.95 ;
        RECT  15.60 7.40 16.30 8.15 ;
        RECT  15.80 3.25 16.30 9.65 ;
        RECT  15.80 8.95 16.65 9.65 ;
    END
END DFRX4
MACRO DLHRSX1
    CLASS CORE ;
    FOREIGN DLHRSX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  10.05 9.30 10.95 10.20 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  19.85 3.70 20.55 8.90 ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  17.15 3.70 17.85 8.90 ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  2.15 6.10 2.65 7.60 ;
        RECT  1.65 6.70 2.65 7.60 ;
        RECT  2.15 6.10 2.85 6.80 ;
        RECT  1.65 6.70 2.85 6.80 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  1.80 10.00 4.55 11.00 ;
        RECT  3.85 9.75 4.55 11.00 ;
        RECT  0.45 10.05 4.55 11.00 ;
        RECT  8.55 7.65 9.25 11.00 ;
        RECT  8.55 7.65 9.45 8.35 ;
        RECT  11.45 7.65 12.15 11.00 ;
        RECT  14.30 7.65 15.00 11.00 ;
        RECT  11.45 10.40 15.00 11.00 ;
        RECT  18.50 7.10 19.20 11.00 ;
        RECT  17.20 10.50 20.55 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.00 2.00 2.70 4.40 ;
        RECT  4.05 2.00 4.75 2.80 ;
        RECT  8.90 2.00 9.60 3.20 ;
        RECT  11.40 2.00 12.15 4.95 ;
        RECT  15.45 2.00 16.15 3.15 ;
        RECT  18.50 2.00 19.20 4.50 ;
        RECT  17.00 2.00 20.55 2.15 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  13.25 3.65 15.05 4.15 ;
        RECT  0.30 2.45 0.80 8.95 ;
        RECT  0.30 2.45 1.00 4.40 ;
        RECT  0.30 7.15 1.15 8.95 ;
        RECT  0.30 3.70 1.35 4.40 ;
        RECT  1.35 4.85 2.05 5.55 ;
        RECT  1.35 4.85 3.85 5.35 ;
        RECT  3.35 3.75 3.85 8.75 ;
        RECT  3.15 7.15 3.85 8.75 ;
        RECT  3.35 3.75 4.05 4.45 ;
        RECT  3.15 8.25 6.45 8.75 ;
        RECT  5.75 8.25 6.45 8.95 ;
        RECT  3.35 3.75 7.45 4.25 ;
        RECT  6.20 9.80 6.90 10.50 ;
        RECT  6.55 2.55 7.25 3.25 ;
        RECT  6.75 3.75 7.45 4.45 ;
        RECT  6.55 2.75 8.40 3.25 ;
        RECT  7.55 6.70 8.05 10.30 ;
        RECT  7.90 2.75 8.05 10.30 ;
        RECT  6.20 9.80 8.05 10.30 ;
        RECT  7.90 2.75 8.40 7.20 ;
        RECT  9.05 4.25 9.80 4.95 ;
        RECT  9.30 6.50 10.00 7.20 ;
        RECT  7.55 6.70 10.00 7.20 ;
        RECT  9.05 4.45 10.95 4.95 ;
        RECT  10.45 4.45 10.95 8.35 ;
        RECT  10.10 7.65 10.95 8.35 ;
        RECT  12.05 6.45 12.75 7.15 ;
        RECT  10.45 6.65 12.75 7.15 ;
        RECT  13.25 3.65 13.75 8.35 ;
        RECT  12.80 7.65 13.75 8.35 ;
        RECT  14.35 2.45 14.45 4.35 ;
        RECT  13.75 2.45 14.45 4.15 ;
        RECT  14.35 3.65 15.05 4.35 ;
        RECT  15.50 3.80 16.35 4.50 ;
        RECT  15.85 3.80 16.35 10.45 ;
        RECT  15.65 7.65 16.35 10.45 ;
        RECT  15.65 9.75 16.75 10.45 ;
    END
END DLHRSX1
MACRO DLHRSX2
    CLASS CORE ;
    FOREIGN DLHRSX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  10.05 9.30 10.95 10.20 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  19.85 2.70 20.55 10.50 ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  17.15 2.70 17.85 10.50 ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  2.15 6.10 2.65 7.60 ;
        RECT  1.65 6.70 2.65 7.60 ;
        RECT  2.15 6.10 2.85 6.80 ;
        RECT  1.65 6.70 2.85 6.80 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  1.80 10.00 4.55 11.00 ;
        RECT  3.85 9.75 4.55 11.00 ;
        RECT  0.45 10.05 4.55 11.00 ;
        RECT  8.55 7.65 9.25 11.00 ;
        RECT  8.55 7.65 9.45 8.35 ;
        RECT  11.45 7.65 12.15 11.00 ;
        RECT  14.30 7.65 15.00 11.00 ;
        RECT  11.45 10.40 15.00 11.00 ;
        RECT  18.50 7.10 19.20 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.00 2.00 2.70 4.40 ;
        RECT  4.05 2.00 4.75 2.80 ;
        RECT  8.90 2.00 9.60 3.20 ;
        RECT  11.40 2.00 12.15 4.95 ;
        RECT  15.45 2.00 16.15 3.15 ;
        RECT  18.50 2.00 19.20 4.50 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  13.25 3.65 15.05 4.15 ;
        RECT  0.30 2.45 0.80 8.95 ;
        RECT  0.30 2.45 1.00 4.40 ;
        RECT  0.30 7.15 1.15 8.95 ;
        RECT  0.30 3.70 1.35 4.40 ;
        RECT  1.35 4.85 2.05 5.55 ;
        RECT  1.35 4.85 3.85 5.35 ;
        RECT  3.35 3.75 3.85 8.75 ;
        RECT  3.15 7.15 3.85 8.75 ;
        RECT  3.35 3.75 4.05 4.45 ;
        RECT  3.15 8.25 6.45 8.75 ;
        RECT  5.75 8.25 6.45 8.95 ;
        RECT  3.35 3.75 7.45 4.25 ;
        RECT  6.20 9.80 6.90 10.50 ;
        RECT  6.55 2.55 7.25 3.25 ;
        RECT  6.75 3.75 7.45 4.45 ;
        RECT  6.55 2.75 8.40 3.25 ;
        RECT  7.55 6.70 8.05 10.30 ;
        RECT  7.90 2.75 8.05 10.30 ;
        RECT  6.20 9.80 8.05 10.30 ;
        RECT  7.90 2.75 8.40 7.20 ;
        RECT  9.05 4.25 9.80 4.95 ;
        RECT  9.30 6.50 10.00 7.20 ;
        RECT  7.55 6.70 10.00 7.20 ;
        RECT  9.05 4.45 10.95 4.95 ;
        RECT  10.45 4.45 10.95 8.35 ;
        RECT  10.10 7.65 10.95 8.35 ;
        RECT  12.05 6.45 12.75 7.15 ;
        RECT  10.45 6.65 12.75 7.15 ;
        RECT  13.25 3.65 13.75 8.35 ;
        RECT  12.80 7.65 13.75 8.35 ;
        RECT  14.35 2.45 14.45 4.35 ;
        RECT  13.75 2.45 14.45 4.15 ;
        RECT  14.35 3.65 15.05 4.35 ;
        RECT  15.50 3.80 16.35 4.50 ;
        RECT  15.85 3.80 16.35 10.45 ;
        RECT  15.65 7.65 16.35 10.45 ;
        RECT  15.65 9.75 16.70 10.45 ;
    END
END DLHRSX2
MACRO DLHRSX4
    CLASS CORE ;
    FOREIGN DLHRSX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  10.05 9.30 10.95 10.20 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  14.25 4.10 15.15 5.00 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  21.30 2.70 22.00 10.50 ;
        RECT  21.25 5.40 22.15 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  18.60 2.70 19.30 10.50 ;
        RECT  18.45 5.40 19.35 6.30 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  2.15 6.10 2.65 7.60 ;
        RECT  1.65 6.70 2.65 7.60 ;
        RECT  2.15 6.10 2.85 6.80 ;
        RECT  1.65 6.70 2.85 6.80 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  1.80 10.00 4.55 11.00 ;
        RECT  3.85 9.75 4.55 11.00 ;
        RECT  0.45 10.05 4.55 11.00 ;
        RECT  8.75 7.65 9.25 11.00 ;
        RECT  8.55 9.75 9.25 11.00 ;
        RECT  8.75 7.65 9.45 8.35 ;
        RECT  11.45 7.65 12.15 11.00 ;
        RECT  14.30 7.65 15.00 11.00 ;
        RECT  17.25 7.10 17.95 11.00 ;
        RECT  19.95 7.10 20.65 11.00 ;
        RECT  22.65 7.10 23.35 11.00 ;
        RECT  0.00 11.00 23.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.00 2.00 2.70 4.40 ;
        RECT  4.05 2.00 4.75 2.80 ;
        RECT  9.10 2.00 9.80 3.25 ;
        RECT  11.45 2.00 12.15 4.95 ;
        RECT  17.25 2.00 17.95 4.50 ;
        RECT  19.95 2.00 20.65 4.50 ;
        RECT  22.65 2.00 23.35 4.50 ;
        RECT  0.00 0.00 23.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.30 2.45 0.80 8.95 ;
        RECT  0.30 2.45 1.00 4.40 ;
        RECT  0.30 7.15 1.15 8.95 ;
        RECT  0.30 3.70 1.35 4.40 ;
        RECT  1.35 4.85 2.05 5.55 ;
        RECT  1.35 4.85 3.85 5.35 ;
        RECT  3.35 3.75 3.85 8.75 ;
        RECT  3.15 7.15 3.85 8.75 ;
        RECT  3.35 3.75 4.05 4.45 ;
        RECT  3.15 8.25 6.45 8.75 ;
        RECT  5.75 8.25 6.45 8.95 ;
        RECT  6.20 9.80 6.90 10.50 ;
        RECT  3.35 3.75 7.70 4.25 ;
        RECT  6.55 2.60 7.25 3.30 ;
        RECT  7.00 3.75 7.70 4.45 ;
        RECT  7.55 6.70 8.05 10.30 ;
        RECT  6.20 9.80 8.05 10.30 ;
        RECT  6.55 2.80 8.65 3.30 ;
        RECT  8.15 2.80 8.65 7.20 ;
        RECT  9.10 4.25 9.85 4.95 ;
        RECT  9.30 6.50 10.00 7.20 ;
        RECT  7.55 6.70 10.00 7.20 ;
        RECT  9.10 4.45 10.95 4.95 ;
        RECT  10.45 4.45 10.95 8.35 ;
        RECT  10.10 7.65 10.95 8.35 ;
        RECT  12.05 6.45 12.75 7.15 ;
        RECT  10.45 6.65 12.75 7.15 ;
        RECT  13.25 2.75 13.75 8.35 ;
        RECT  12.80 7.65 13.75 8.35 ;
        RECT  13.25 5.50 15.35 6.00 ;
        RECT  13.95 2.55 14.65 3.25 ;
        RECT  13.25 2.75 14.65 3.25 ;
        RECT  14.65 5.50 15.35 6.20 ;
        RECT  15.85 3.75 16.35 10.45 ;
        RECT  15.65 7.65 16.35 10.45 ;
        RECT  15.75 3.75 16.45 4.45 ;
        RECT  15.65 9.75 16.70 10.45 ;
    END
END DLHRSX4
MACRO DLHRX1
    CLASS CORE ;
    FOREIGN DLHRX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.35 15.15 6.35 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  17.15 3.75 17.95 4.45 ;
        RECT  17.05 5.35 17.95 6.35 ;
        RECT  17.35 3.75 17.95 8.90 ;
        RECT  17.15 7.15 17.95 8.90 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  19.85 3.75 20.35 8.90 ;
        RECT  19.85 3.75 20.55 4.45 ;
        RECT  19.85 7.15 20.55 8.90 ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  2.15 6.10 2.65 7.60 ;
        RECT  1.65 6.70 2.65 7.60 ;
        RECT  2.15 6.10 2.85 6.80 ;
        RECT  1.65 6.70 2.85 6.80 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.30 5.40 5.35 6.30 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  1.80 10.00 4.55 11.00 ;
        RECT  3.85 9.75 4.55 11.00 ;
        RECT  0.45 10.05 4.55 11.00 ;
        RECT  8.70 7.75 9.40 11.00 ;
        RECT  14.30 7.60 15.00 11.00 ;
        RECT  18.50 7.15 19.20 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.00 2.00 2.70 4.40 ;
        RECT  3.70 2.00 4.40 2.80 ;
        RECT  8.70 2.00 9.40 3.25 ;
        RECT  11.45 2.00 12.15 3.25 ;
        RECT  14.30 2.00 15.00 3.65 ;
        RECT  18.50 2.00 19.20 4.45 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.30 2.45 0.80 8.95 ;
        RECT  0.30 2.45 1.00 4.40 ;
        RECT  0.30 7.15 1.15 8.95 ;
        RECT  0.30 3.70 1.35 4.40 ;
        RECT  1.35 4.85 2.05 5.55 ;
        RECT  1.35 4.85 3.85 5.35 ;
        RECT  3.35 3.75 3.85 8.90 ;
        RECT  3.15 7.15 3.85 8.90 ;
        RECT  3.35 3.75 4.05 4.45 ;
        RECT  3.15 8.40 6.45 8.90 ;
        RECT  5.75 8.40 6.45 9.10 ;
        RECT  6.20 2.55 6.90 3.25 ;
        RECT  6.20 9.75 6.90 10.45 ;
        RECT  6.55 3.75 7.25 4.45 ;
        RECT  3.35 3.95 7.25 4.45 ;
        RECT  6.20 2.75 8.25 3.25 ;
        RECT  7.55 6.65 8.05 10.25 ;
        RECT  7.75 2.75 8.05 10.25 ;
        RECT  6.20 9.75 8.05 10.25 ;
        RECT  7.75 2.75 8.25 7.15 ;
        RECT  9.15 3.75 9.85 4.45 ;
        RECT  7.75 3.95 9.85 4.45 ;
        RECT  10.05 2.55 10.95 3.25 ;
        RECT  10.45 2.55 10.95 4.25 ;
        RECT  10.40 6.45 11.10 7.15 ;
        RECT  7.55 6.65 11.10 7.15 ;
        RECT  10.45 3.75 12.45 4.25 ;
        RECT  11.05 7.75 11.75 10.50 ;
        RECT  11.75 3.75 12.25 8.30 ;
        RECT  11.05 7.75 12.25 8.30 ;
        RECT  11.75 3.75 12.45 4.45 ;
        RECT  11.75 6.45 12.45 7.15 ;
        RECT  12.95 2.55 13.45 10.50 ;
        RECT  12.80 2.55 13.50 3.25 ;
        RECT  12.95 7.60 13.65 10.50 ;
        RECT  12.60 9.80 13.65 10.50 ;
        RECT  13.95 4.15 14.65 4.85 ;
        RECT  15.65 2.95 16.35 3.65 ;
        RECT  13.95 4.35 16.35 4.85 ;
        RECT  15.85 2.95 16.35 9.40 ;
        RECT  15.65 7.60 16.35 9.40 ;
    END
END DLHRX1
MACRO DLHRX2
    CLASS CORE ;
    FOREIGN DLHRX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.35 15.15 6.35 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  17.15 2.70 17.95 4.50 ;
        RECT  17.05 5.35 17.95 6.35 ;
        RECT  17.35 2.70 17.95 10.55 ;
        RECT  17.15 7.15 17.95 10.55 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  19.85 2.70 20.35 10.55 ;
        RECT  19.85 2.70 20.55 4.50 ;
        RECT  19.85 7.15 20.55 10.55 ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  2.15 6.10 2.65 7.60 ;
        RECT  1.65 6.70 2.65 7.60 ;
        RECT  2.15 6.10 2.85 6.80 ;
        RECT  1.65 6.70 2.85 6.80 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.30 5.40 5.35 6.30 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  1.80 10.00 4.55 11.00 ;
        RECT  3.85 9.75 4.55 11.00 ;
        RECT  0.45 10.05 4.55 11.00 ;
        RECT  8.70 7.75 9.40 11.00 ;
        RECT  14.30 7.60 15.00 11.00 ;
        RECT  18.50 7.15 19.20 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.00 2.00 2.70 4.40 ;
        RECT  3.70 2.00 4.40 2.80 ;
        RECT  8.70 2.00 9.40 3.25 ;
        RECT  11.45 2.00 12.15 3.25 ;
        RECT  14.30 2.00 15.00 3.65 ;
        RECT  18.50 2.00 19.20 4.50 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.30 2.45 0.80 8.95 ;
        RECT  0.30 2.45 1.00 4.40 ;
        RECT  0.30 7.15 1.15 8.95 ;
        RECT  0.30 3.70 1.35 4.40 ;
        RECT  1.35 4.85 2.05 5.55 ;
        RECT  1.35 4.85 3.85 5.35 ;
        RECT  3.35 3.75 3.85 8.90 ;
        RECT  3.15 7.15 3.85 8.90 ;
        RECT  3.35 3.75 4.05 4.45 ;
        RECT  3.15 8.40 6.45 8.90 ;
        RECT  5.75 8.40 6.45 9.10 ;
        RECT  6.20 2.55 6.90 3.25 ;
        RECT  6.20 9.75 6.90 10.45 ;
        RECT  6.55 3.75 7.25 4.45 ;
        RECT  3.35 3.95 7.25 4.45 ;
        RECT  6.20 2.75 8.25 3.25 ;
        RECT  7.55 6.65 8.05 10.25 ;
        RECT  7.75 2.75 8.05 10.25 ;
        RECT  6.20 9.75 8.05 10.25 ;
        RECT  7.75 2.75 8.25 7.15 ;
        RECT  9.15 3.75 9.85 4.45 ;
        RECT  7.75 3.95 9.85 4.45 ;
        RECT  10.05 2.55 10.95 3.25 ;
        RECT  10.45 2.55 10.95 4.25 ;
        RECT  10.40 6.45 11.10 7.15 ;
        RECT  7.55 6.65 11.10 7.15 ;
        RECT  10.45 3.75 12.45 4.25 ;
        RECT  11.05 7.75 11.75 10.50 ;
        RECT  11.75 3.75 12.25 8.30 ;
        RECT  11.05 7.75 12.25 8.30 ;
        RECT  11.75 3.75 12.45 4.45 ;
        RECT  11.75 6.45 12.45 7.15 ;
        RECT  12.95 2.55 13.45 10.50 ;
        RECT  12.80 2.55 13.50 3.25 ;
        RECT  12.95 7.60 13.65 10.50 ;
        RECT  12.60 9.80 13.65 10.50 ;
        RECT  13.95 4.15 14.65 4.85 ;
        RECT  15.65 2.95 16.35 3.65 ;
        RECT  13.95 4.35 16.35 4.85 ;
        RECT  15.85 2.95 16.35 9.40 ;
        RECT  15.65 7.60 16.35 9.40 ;
    END
END DLHRX2
MACRO DLHRX4
    CLASS CORE ;
    FOREIGN DLHRX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.35 15.15 6.35 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.40 19.35 6.30 ;
        RECT  18.55 2.70 19.35 10.55 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  21.25 2.70 21.95 10.55 ;
        RECT  21.25 5.40 22.15 6.30 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  2.15 6.10 2.65 7.60 ;
        RECT  1.65 6.70 2.65 7.60 ;
        RECT  2.15 6.10 2.85 6.80 ;
        RECT  1.65 6.70 2.85 6.80 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.30 5.40 5.35 6.30 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  1.80 10.00 4.55 11.00 ;
        RECT  3.85 9.75 4.55 11.00 ;
        RECT  0.45 10.05 4.55 11.00 ;
        RECT  8.70 7.75 9.40 11.00 ;
        RECT  14.30 7.60 15.00 11.00 ;
        RECT  17.20 7.15 17.90 11.00 ;
        RECT  19.90 7.15 20.60 11.00 ;
        RECT  22.60 7.15 23.30 11.00 ;
        RECT  0.00 11.00 23.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.00 2.00 2.70 4.40 ;
        RECT  3.70 2.00 4.40 2.80 ;
        RECT  8.70 2.00 9.40 3.25 ;
        RECT  11.45 2.00 12.15 3.25 ;
        RECT  14.30 2.00 15.00 3.65 ;
        RECT  17.20 2.00 17.90 4.50 ;
        RECT  19.90 2.00 20.60 4.50 ;
        RECT  22.60 2.00 23.30 4.50 ;
        RECT  0.00 0.00 23.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.30 2.45 0.80 8.95 ;
        RECT  0.30 2.45 1.00 4.40 ;
        RECT  0.30 7.15 1.15 8.95 ;
        RECT  0.30 3.70 1.35 4.40 ;
        RECT  1.35 4.85 2.05 5.55 ;
        RECT  1.35 4.85 3.85 5.35 ;
        RECT  3.35 3.75 3.85 8.90 ;
        RECT  3.15 7.15 3.85 8.90 ;
        RECT  3.35 3.75 4.05 4.45 ;
        RECT  3.15 8.40 6.45 8.90 ;
        RECT  5.75 8.40 6.45 9.10 ;
        RECT  6.20 2.55 6.90 3.25 ;
        RECT  6.20 9.75 6.90 10.45 ;
        RECT  6.55 3.75 7.25 4.45 ;
        RECT  3.35 3.95 7.25 4.45 ;
        RECT  6.20 2.75 8.25 3.25 ;
        RECT  7.55 6.65 8.05 10.25 ;
        RECT  7.75 2.75 8.05 10.25 ;
        RECT  6.20 9.75 8.05 10.25 ;
        RECT  7.75 2.75 8.25 7.15 ;
        RECT  9.15 3.75 9.85 4.45 ;
        RECT  7.75 3.95 9.85 4.45 ;
        RECT  10.05 2.55 10.95 3.25 ;
        RECT  10.45 2.55 10.95 4.25 ;
        RECT  10.40 6.45 11.10 7.15 ;
        RECT  7.55 6.65 11.10 7.15 ;
        RECT  10.45 3.75 12.45 4.25 ;
        RECT  11.05 7.75 11.75 10.50 ;
        RECT  11.75 3.75 12.25 8.30 ;
        RECT  11.05 7.75 12.25 8.30 ;
        RECT  11.75 3.75 12.45 4.45 ;
        RECT  11.75 6.45 12.45 7.15 ;
        RECT  12.95 2.55 13.45 10.50 ;
        RECT  12.80 2.55 13.50 3.25 ;
        RECT  12.95 7.60 13.65 10.50 ;
        RECT  12.60 9.80 13.65 10.50 ;
        RECT  13.95 4.15 14.65 4.85 ;
        RECT  15.65 2.95 16.35 3.65 ;
        RECT  13.95 4.35 16.35 4.85 ;
        RECT  15.85 2.95 16.35 9.40 ;
        RECT  15.65 7.60 16.35 9.40 ;
    END
END DLHRX4
MACRO DLHSX1
    CLASS CORE ;
    FOREIGN DLHSX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.55 5.00 ;
        RECT  8.65 4.10 9.70 4.80 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  17.05 3.75 17.75 9.65 ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  14.35 3.75 15.05 9.65 ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  2.15 6.10 2.65 7.60 ;
        RECT  1.65 6.70 2.65 7.60 ;
        RECT  2.15 6.10 2.85 6.80 ;
        RECT  1.65 6.70 2.85 6.80 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.30 5.40 5.35 6.30 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  1.80 10.00 4.55 11.00 ;
        RECT  3.85 9.75 4.55 11.00 ;
        RECT  0.45 10.05 4.55 11.00 ;
        RECT  8.20 7.35 9.05 8.05 ;
        RECT  8.55 7.35 9.05 11.00 ;
        RECT  8.55 8.60 9.25 11.00 ;
        RECT  11.05 7.40 11.75 9.10 ;
        RECT  8.55 8.60 11.75 9.10 ;
        RECT  15.70 7.90 16.40 11.00 ;
        RECT  10.05 10.55 17.75 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.00 2.00 2.70 4.40 ;
        RECT  3.70 2.00 4.40 2.80 ;
        RECT  8.55 2.00 9.25 3.60 ;
        RECT  12.65 2.00 13.35 3.15 ;
        RECT  15.70 2.00 16.40 4.45 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.30 2.45 0.80 8.95 ;
        RECT  0.30 2.45 1.00 4.40 ;
        RECT  0.30 7.15 1.15 8.95 ;
        RECT  0.30 3.70 1.35 4.40 ;
        RECT  1.35 4.85 2.05 5.55 ;
        RECT  1.35 4.85 3.85 5.35 ;
        RECT  3.35 3.75 3.85 8.90 ;
        RECT  3.15 7.15 3.85 8.90 ;
        RECT  3.35 3.75 4.05 4.90 ;
        RECT  3.15 8.40 6.25 8.90 ;
        RECT  5.55 8.40 6.25 9.10 ;
        RECT  3.35 4.40 7.10 4.90 ;
        RECT  6.20 2.95 6.90 3.65 ;
        RECT  6.20 9.75 6.90 10.45 ;
        RECT  6.40 4.20 7.10 4.90 ;
        RECT  1.35 4.85 7.10 4.90 ;
        RECT  6.20 3.15 8.05 3.65 ;
        RECT  7.25 5.50 7.75 10.25 ;
        RECT  7.55 3.15 7.75 10.25 ;
        RECT  6.20 9.75 7.75 10.25 ;
        RECT  7.55 3.15 8.05 6.00 ;
        RECT  9.55 6.45 10.25 8.05 ;
        RECT  10.15 5.30 10.85 6.00 ;
        RECT  7.25 5.50 10.85 6.00 ;
        RECT  10.90 2.95 11.90 3.65 ;
        RECT  11.40 2.95 11.90 6.95 ;
        RECT  11.40 6.25 12.10 6.95 ;
        RECT  9.55 6.45 12.10 6.95 ;
        RECT  12.70 3.80 13.40 4.50 ;
        RECT  12.90 3.80 13.10 9.10 ;
        RECT  12.40 7.30 13.10 9.10 ;
        RECT  12.90 3.80 13.40 7.80 ;
        RECT  12.40 7.30 13.40 7.80 ;
        RECT  12.90 6.25 13.60 6.95 ;
    END
END DLHSX1
MACRO DLHSX2
    CLASS CORE ;
    FOREIGN DLHSX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.55 5.00 ;
        RECT  8.65 4.10 9.70 4.80 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  17.05 2.75 17.75 10.55 ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  14.35 2.75 15.05 10.55 ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  2.15 6.10 2.65 7.60 ;
        RECT  1.65 6.70 2.65 7.60 ;
        RECT  2.15 6.10 2.85 6.80 ;
        RECT  1.65 6.70 2.85 6.80 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.30 5.40 5.35 6.30 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  1.80 10.00 4.55 11.00 ;
        RECT  3.85 9.75 4.55 11.00 ;
        RECT  0.45 10.05 4.55 11.00 ;
        RECT  8.20 7.35 9.05 8.05 ;
        RECT  8.55 7.35 9.05 11.00 ;
        RECT  8.55 8.60 9.25 11.00 ;
        RECT  11.05 7.40 11.75 9.10 ;
        RECT  8.55 8.60 11.75 9.10 ;
        RECT  10.05 10.55 13.55 11.00 ;
        RECT  15.70 7.10 16.40 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.00 2.00 2.70 4.40 ;
        RECT  3.70 2.00 4.40 2.80 ;
        RECT  8.55 2.00 9.25 3.60 ;
        RECT  12.65 2.00 13.35 3.15 ;
        RECT  15.70 2.00 16.40 4.45 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.30 2.45 0.80 8.95 ;
        RECT  0.30 2.45 1.00 4.40 ;
        RECT  0.30 7.15 1.15 8.95 ;
        RECT  0.30 3.70 1.35 4.40 ;
        RECT  1.35 4.85 2.05 5.55 ;
        RECT  1.35 4.85 3.85 5.35 ;
        RECT  3.35 3.75 3.85 8.90 ;
        RECT  3.15 7.15 3.85 8.90 ;
        RECT  3.35 3.75 4.05 4.90 ;
        RECT  3.15 8.40 6.25 8.90 ;
        RECT  5.55 8.40 6.25 9.10 ;
        RECT  3.35 4.40 7.10 4.90 ;
        RECT  6.20 2.95 6.90 3.65 ;
        RECT  6.20 9.75 6.90 10.45 ;
        RECT  6.40 4.20 7.10 4.90 ;
        RECT  1.35 4.85 7.10 4.90 ;
        RECT  6.20 3.15 8.05 3.65 ;
        RECT  7.25 5.50 7.75 10.25 ;
        RECT  7.55 3.15 7.75 10.25 ;
        RECT  6.20 9.75 7.75 10.25 ;
        RECT  7.55 3.15 8.05 6.00 ;
        RECT  9.55 6.45 10.25 8.05 ;
        RECT  10.15 5.30 10.85 6.00 ;
        RECT  7.25 5.50 10.85 6.00 ;
        RECT  10.90 2.95 11.90 3.65 ;
        RECT  11.40 2.95 11.90 6.95 ;
        RECT  11.40 6.25 12.10 6.95 ;
        RECT  9.55 6.45 12.10 6.95 ;
        RECT  12.70 3.80 13.40 4.50 ;
        RECT  12.90 3.80 13.10 9.10 ;
        RECT  12.40 7.30 13.10 9.10 ;
        RECT  12.90 3.80 13.40 7.80 ;
        RECT  12.40 7.30 13.40 7.80 ;
        RECT  12.90 6.25 13.60 6.95 ;
    END
END DLHSX2
MACRO DLHSX4
    CLASS CORE ;
    FOREIGN DLHSX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.55 5.00 ;
        RECT  8.65 4.10 9.70 4.80 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  18.45 2.75 19.15 10.55 ;
        RECT  18.45 5.40 19.35 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  15.75 2.75 16.45 10.55 ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  2.15 6.10 2.65 7.60 ;
        RECT  1.65 6.70 2.65 7.60 ;
        RECT  2.15 6.10 2.85 6.80 ;
        RECT  1.65 6.70 2.85 6.80 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.30 5.40 5.35 6.30 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  1.80 10.00 4.55 11.00 ;
        RECT  3.85 9.75 4.55 11.00 ;
        RECT  0.45 10.05 4.55 11.00 ;
        RECT  8.20 7.35 9.05 8.05 ;
        RECT  8.55 7.35 9.05 11.00 ;
        RECT  8.55 8.60 9.25 11.00 ;
        RECT  11.05 7.40 11.75 9.10 ;
        RECT  8.55 8.60 11.75 9.10 ;
        RECT  10.05 10.55 13.55 11.00 ;
        RECT  14.40 7.10 15.10 11.00 ;
        RECT  17.10 7.10 17.80 11.00 ;
        RECT  19.80 7.10 20.50 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.00 2.00 2.70 4.40 ;
        RECT  3.70 2.00 4.40 2.80 ;
        RECT  8.55 2.00 9.25 3.60 ;
        RECT  12.65 2.00 13.35 3.15 ;
        RECT  14.40 2.00 15.10 4.45 ;
        RECT  17.10 2.00 17.80 4.45 ;
        RECT  19.80 2.00 20.50 4.45 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.30 2.45 0.80 8.95 ;
        RECT  0.30 2.45 1.00 4.40 ;
        RECT  0.30 7.15 1.15 8.95 ;
        RECT  0.30 3.70 1.35 4.40 ;
        RECT  1.35 4.85 2.05 5.55 ;
        RECT  1.35 4.85 3.85 5.35 ;
        RECT  3.35 3.75 3.85 8.90 ;
        RECT  3.15 7.15 3.85 8.90 ;
        RECT  3.35 3.75 4.05 4.90 ;
        RECT  3.15 8.40 6.25 8.90 ;
        RECT  5.55 8.40 6.25 9.10 ;
        RECT  3.35 4.40 7.10 4.90 ;
        RECT  6.20 2.95 6.90 3.65 ;
        RECT  6.20 9.75 6.90 10.45 ;
        RECT  6.40 4.20 7.10 4.90 ;
        RECT  1.35 4.85 7.10 4.90 ;
        RECT  6.20 3.15 8.05 3.65 ;
        RECT  7.25 5.50 7.75 10.25 ;
        RECT  7.55 3.15 7.75 10.25 ;
        RECT  6.20 9.75 7.75 10.25 ;
        RECT  7.55 3.15 8.05 6.00 ;
        RECT  9.55 6.45 10.25 8.05 ;
        RECT  10.15 5.30 10.85 6.00 ;
        RECT  7.25 5.50 10.85 6.00 ;
        RECT  10.90 2.95 11.90 3.65 ;
        RECT  11.40 2.95 11.90 6.95 ;
        RECT  11.40 6.25 12.10 6.95 ;
        RECT  9.55 6.45 12.10 6.95 ;
        RECT  12.70 3.80 13.40 4.50 ;
        RECT  12.90 3.80 13.10 9.10 ;
        RECT  12.40 7.30 13.10 9.10 ;
        RECT  12.90 3.80 13.40 7.80 ;
        RECT  12.40 7.30 13.40 7.80 ;
        RECT  12.90 6.25 13.60 6.95 ;
    END
END DLHSX4
#MACRO DLHX1
#    CLASS CORE ;
#    FOREIGN DLHX1 0.00 0.00  ;
#    ORIGIN 0.00 0.00 ;
#    SIZE 15.40 BY 13.00 ;
#    SYMMETRY x y r90 ;
#    SITE core ;
#    PIN QN
#        DIRECTION OUTPUT ;
#        ANTENNADIFFAREA 1.0 ;
#        PORT
#        LAYER M1M ;
#        RECT  14.25 3.75 14.95 8.90 ;
#        RECT  14.25 5.40 15.15 6.30 ;
#        END
#    END QN
#    PIN Q
#        DIRECTION OUTPUT ;
#        ANTENNADIFFAREA 1.0 ;
#        PORT
#        LAYER M1M ;
#        RECT  11.55 3.75 12.25 8.90 ;
#        RECT  11.45 5.40 12.35 6.30 ;
#        END
#    END Q
#    PIN G
#        DIRECTION INPUT ;
#        ANTENNAGATEAREA 1.05 ;
#        PORT
#        LAYER M1M ;
#        RECT  2.15 6.10 2.65 7.60 ;
#        RECT  1.65 6.70 2.65 7.60 ;
#        RECT  2.15 6.10 2.85 6.80 ;
#        RECT  1.65 6.70 2.85 6.80 ;
#        END
#    END G
#    PIN D
#        DIRECTION INPUT ;
#        ANTENNAGATEAREA 1.05 ;
#        PORT
#        LAYER M1M ;
#        RECT  4.40 6.70 5.35 7.75 ;
#        END
#    END D
#    PIN vdd!
#        DIRECTION INOUT ;
#        USE power ;
#        SHAPE ABUTMENT ;
#        PORT
#        LAYER M1M ;
#        RECT  1.80 8.10 2.50 11.00 ;
#        RECT  1.80 9.75 4.20 11.00 ;
#        RECT  0.45 10.05 4.20 11.00 ;
#        RECT  8.70 7.10 9.40 11.00 ;
#        RECT  12.90 7.15 13.60 11.00 ;
#        RECT  7.50 10.05 14.95 11.00 ;
#        RECT  0.00 11.00 15.40 13.00 ;
#        END
#    END vdd!
#    PIN gnd!
#        DIRECTION INOUT ;
#        USE ground ;
#        SHAPE ABUTMENT ;
#        PORT
#        LAYER M1M ;
#        RECT  2.00 2.00 2.70 4.40 ;
#        RECT  3.70 2.00 4.40 2.80 ;
#        RECT  8.70 2.00 9.40 4.50 ;
#        RECT  12.90 2.00 13.60 4.45 ;
#        RECT  0.00 0.00 15.40 2.00 ;
#        END
#    END gnd!
#    OBS
#        LAYER M1M ;
#        RECT  0.30 2.45 0.80 8.95 ;
#        RECT  0.30 2.45 1.00 4.40 ;
#        RECT  0.30 7.15 1.15 8.95 ;
#        RECT  0.30 3.70 1.35 4.40 ;
#        RECT  1.35 4.85 2.05 5.55 ;
#        RECT  1.35 4.85 4.05 5.35 ;
#        RECT  3.35 3.75 3.85 8.90 ;
#        RECT  3.15 7.15 3.85 8.90 ;
#        RECT  3.35 3.75 4.05 5.90 ;
#        RECT  3.15 8.40 5.90 8.90 ;
#        RECT  5.20 8.40 5.90 9.10 ;
#        RECT  6.20 2.50 6.90 4.50 ;
#        RECT  6.35 7.10 7.05 10.45 ;
#        RECT  5.85 9.75 7.05 10.45 ;
#        RECT  6.40 5.20 7.10 5.90 ;
#        RECT  3.35 5.40 7.10 5.90 ;
#        RECT  6.20 4.00 8.05 4.50 ;
#        RECT  7.55 4.00 8.05 7.80 ;
#        RECT  6.35 7.10 8.05 7.80 ;
#        RECT  9.10 5.80 9.80 6.50 ;
#        RECT  7.55 6.00 9.80 6.50 ;
#        RECT  10.05 2.65 10.75 4.50 ;
#        RECT  10.25 2.65 10.75 8.90 ;
#        RECT  10.05 7.10 10.75 8.90 ;
#        RECT  10.05 2.65 11.10 3.35 ;
#    END
#END DLHX1
MACRO DLHX2
    CLASS CORE ;
    FOREIGN DLHX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  14.25 2.70 14.95 10.55 ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.55 2.70 12.25 10.55 ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  2.15 6.10 2.65 7.60 ;
        RECT  1.65 6.70 2.65 7.60 ;
        RECT  2.15 6.10 2.85 6.80 ;
        RECT  1.65 6.70 2.85 6.80 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.40 6.70 5.35 7.75 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  1.80 9.75 4.20 11.00 ;
        RECT  0.45 10.05 4.20 11.00 ;
        RECT  8.70 7.10 9.40 11.00 ;
        RECT  7.50 10.05 10.75 11.00 ;
        RECT  12.90 7.10 13.60 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.00 2.00 2.70 4.40 ;
        RECT  3.70 2.00 4.40 2.80 ;
        RECT  8.70 2.00 9.40 4.50 ;
        RECT  12.90 2.00 13.60 4.45 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.30 2.45 0.80 8.95 ;
        RECT  0.30 2.45 1.00 4.40 ;
        RECT  0.30 7.15 1.15 8.95 ;
        RECT  0.30 3.70 1.35 4.40 ;
        RECT  1.35 4.85 2.05 5.55 ;
        RECT  1.35 4.85 4.05 5.35 ;
        RECT  3.35 3.75 3.85 8.90 ;
        RECT  3.15 7.15 3.85 8.90 ;
        RECT  3.35 3.75 4.05 5.90 ;
        RECT  3.15 8.40 5.90 8.90 ;
        RECT  5.20 8.40 5.90 9.10 ;
        RECT  6.20 2.50 6.90 4.50 ;
        RECT  6.35 7.10 7.05 10.45 ;
        RECT  5.85 9.75 7.05 10.45 ;
        RECT  6.40 5.20 7.10 5.90 ;
        RECT  3.35 5.40 7.10 5.90 ;
        RECT  6.20 4.00 8.05 4.50 ;
        RECT  7.55 4.00 8.05 7.80 ;
        RECT  6.35 7.10 8.05 7.80 ;
        RECT  9.10 5.80 9.80 6.50 ;
        RECT  7.55 6.00 9.80 6.50 ;
        RECT  10.05 2.65 10.75 4.50 ;
        RECT  10.25 2.65 10.75 8.90 ;
        RECT  10.05 7.10 10.75 8.90 ;
        RECT  10.05 2.65 11.10 3.35 ;
    END
END DLHX2
MACRO DLHX4
    CLASS CORE ;
    FOREIGN DLHX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  15.65 2.70 16.35 10.55 ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  12.95 2.70 13.65 10.55 ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  2.15 6.10 2.65 7.60 ;
        RECT  1.65 6.70 2.65 7.60 ;
        RECT  2.15 6.10 2.85 6.80 ;
        RECT  1.65 6.70 2.85 6.80 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.40 6.70 5.35 7.75 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  1.80 9.75 4.20 11.00 ;
        RECT  0.45 10.05 4.20 11.00 ;
        RECT  8.70 7.10 9.40 11.00 ;
        RECT  7.50 10.05 10.75 11.00 ;
        RECT  11.60 7.10 12.30 11.00 ;
        RECT  14.30 7.10 15.00 11.00 ;
        RECT  17.00 7.10 17.70 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.00 2.00 2.70 4.40 ;
        RECT  3.70 2.00 4.40 2.80 ;
        RECT  8.70 2.00 9.40 4.50 ;
        RECT  11.60 2.00 12.30 4.45 ;
        RECT  14.30 2.00 15.00 4.45 ;
        RECT  17.00 2.00 17.70 4.45 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.30 2.45 0.80 8.95 ;
        RECT  0.30 2.45 1.00 4.40 ;
        RECT  0.30 7.15 1.15 8.95 ;
        RECT  0.30 3.70 1.35 4.40 ;
        RECT  1.35 4.85 2.05 5.55 ;
        RECT  1.35 4.85 4.05 5.35 ;
        RECT  3.35 3.75 3.85 8.90 ;
        RECT  3.15 7.15 3.85 8.90 ;
        RECT  3.35 3.75 4.05 5.90 ;
        RECT  3.15 8.40 5.90 8.90 ;
        RECT  5.20 8.40 5.90 9.10 ;
        RECT  6.20 2.50 6.90 4.50 ;
        RECT  6.35 7.10 7.05 10.45 ;
        RECT  5.85 9.75 7.05 10.45 ;
        RECT  6.40 5.20 7.10 5.90 ;
        RECT  3.35 5.40 7.10 5.90 ;
        RECT  6.20 4.00 8.05 4.50 ;
        RECT  7.55 4.00 8.05 7.80 ;
        RECT  6.35 7.10 8.05 7.80 ;
        RECT  9.10 5.80 9.80 6.50 ;
        RECT  7.55 6.00 9.80 6.50 ;
        RECT  10.05 2.65 10.75 4.50 ;
        RECT  10.25 2.65 10.75 8.90 ;
        RECT  10.05 7.10 10.75 8.90 ;
        RECT  10.05 2.65 11.10 3.35 ;
    END
END DLHX4
MACRO DLLRSX1
    CLASS CORE ;
    FOREIGN DLLRSX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  10.05 9.30 10.95 10.20 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  14.25 3.75 14.95 5.00 ;
        RECT  14.25 4.00 15.15 5.00 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  19.85 2.50 20.55 3.20 ;
        RECT  20.05 2.50 20.55 9.35 ;
        RECT  19.85 7.60 20.55 9.35 ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  17.15 2.50 17.35 9.35 ;
        RECT  16.85 2.50 17.35 6.30 ;
        RECT  17.15 5.40 17.65 9.35 ;
        RECT  17.15 7.60 17.85 9.35 ;
        RECT  16.85 2.50 17.95 3.20 ;
        RECT  16.85 5.40 17.95 6.30 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.60 5.35 2.60 6.35 ;
        RECT  1.25 5.65 2.60 6.35 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.30 4.25 6.80 4.95 ;
        RECT  5.80 4.05 6.80 5.05 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.15 2.50 11.00 ;
        RECT  3.85 9.70 4.55 11.00 ;
        RECT  0.45 10.05 4.55 11.00 ;
        RECT  8.75 7.65 9.25 11.00 ;
        RECT  8.55 9.70 9.25 11.00 ;
        RECT  8.75 7.65 9.45 8.35 ;
        RECT  11.45 7.65 12.15 11.00 ;
        RECT  14.30 7.65 15.00 11.00 ;
        RECT  18.50 7.60 19.20 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.35 ;
        RECT  3.85 2.00 4.55 3.25 ;
        RECT  8.75 2.00 9.45 3.25 ;
        RECT  11.75 2.00 12.50 4.95 ;
        RECT  11.55 4.20 12.50 4.95 ;
        RECT  18.50 2.00 19.20 4.85 ;
        RECT  17.85 4.15 19.20 4.85 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.50 3.70 3.65 4.20 ;
        RECT  0.25 4.35 0.75 8.85 ;
        RECT  0.25 7.15 1.15 8.85 ;
        RECT  1.00 3.10 1.80 4.85 ;
        RECT  0.25 4.35 1.80 4.85 ;
        RECT  3.15 2.55 3.20 8.90 ;
        RECT  2.50 2.55 3.20 4.20 ;
        RECT  3.15 3.70 3.65 8.90 ;
        RECT  3.15 7.15 3.85 8.90 ;
        RECT  3.15 8.40 6.45 8.90 ;
        RECT  5.75 8.40 6.45 9.10 ;
        RECT  3.15 5.55 7.25 6.05 ;
        RECT  6.20 2.55 6.90 3.25 ;
        RECT  6.20 9.75 6.90 10.45 ;
        RECT  6.55 5.55 7.25 6.25 ;
        RECT  6.20 2.75 8.25 3.25 ;
        RECT  7.55 6.65 8.05 10.25 ;
        RECT  7.75 2.75 8.05 10.25 ;
        RECT  6.20 9.75 8.05 10.25 ;
        RECT  7.75 2.75 8.25 7.15 ;
        RECT  9.10 4.25 9.85 4.95 ;
        RECT  9.25 6.45 9.95 7.15 ;
        RECT  7.55 6.65 9.95 7.15 ;
        RECT  9.10 4.45 10.95 4.95 ;
        RECT  10.45 4.45 10.95 8.35 ;
        RECT  10.10 7.65 10.95 8.35 ;
        RECT  12.05 6.45 12.75 7.15 ;
        RECT  10.45 6.65 12.75 7.15 ;
        RECT  13.25 2.75 13.75 8.35 ;
        RECT  12.80 7.65 13.75 8.35 ;
        RECT  13.25 5.50 15.35 6.00 ;
        RECT  14.15 2.55 14.85 3.25 ;
        RECT  13.25 2.75 14.85 3.25 ;
        RECT  14.65 5.50 15.35 6.20 ;
        RECT  15.65 3.10 16.35 4.95 ;
        RECT  15.85 3.10 16.35 9.40 ;
        RECT  15.65 7.65 16.35 9.40 ;
    END
END DLLRSX1
MACRO DLLRSX2
    CLASS CORE ;
    FOREIGN DLLRSX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  10.05 9.30 10.95 10.20 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  14.25 3.75 14.95 5.00 ;
        RECT  14.25 4.00 15.15 5.00 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  19.85 2.50 20.55 3.20 ;
        RECT  20.05 2.50 20.55 10.50 ;
        RECT  19.85 7.60 20.55 10.50 ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  17.15 2.50 17.35 10.50 ;
        RECT  16.85 2.50 17.35 6.30 ;
        RECT  17.15 5.40 17.65 10.50 ;
        RECT  17.15 7.60 17.85 10.50 ;
        RECT  16.85 2.50 17.95 3.20 ;
        RECT  16.85 5.40 17.95 6.30 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.60 5.35 2.60 6.35 ;
        RECT  1.25 5.65 2.60 6.35 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.30 4.25 6.80 4.95 ;
        RECT  5.80 4.05 6.80 5.05 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.15 2.50 11.00 ;
        RECT  3.85 9.70 4.55 11.00 ;
        RECT  0.45 10.05 4.55 11.00 ;
        RECT  8.70 7.65 9.25 11.00 ;
        RECT  8.55 9.70 9.25 11.00 ;
        RECT  8.70 7.65 9.40 8.35 ;
        RECT  11.40 7.65 12.10 8.35 ;
        RECT  11.50 7.65 12.10 11.00 ;
        RECT  14.25 7.65 14.95 11.00 ;
        RECT  18.50 7.60 19.20 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.35 ;
        RECT  3.85 2.00 4.55 3.25 ;
        RECT  8.75 2.00 9.45 3.25 ;
        RECT  11.75 2.00 12.45 4.95 ;
        RECT  11.40 4.20 12.45 4.95 ;
        RECT  18.50 2.00 19.20 4.85 ;
        RECT  17.85 4.15 19.20 4.85 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.50 3.70 3.65 4.20 ;
        RECT  0.25 4.35 0.75 8.85 ;
        RECT  0.25 7.15 1.15 8.85 ;
        RECT  1.00 3.10 1.80 4.85 ;
        RECT  0.25 4.35 1.80 4.85 ;
        RECT  3.15 2.55 3.20 8.90 ;
        RECT  2.50 2.55 3.20 4.20 ;
        RECT  3.15 3.70 3.65 8.90 ;
        RECT  3.15 7.15 3.85 8.90 ;
        RECT  3.15 8.40 6.45 8.90 ;
        RECT  5.75 8.40 6.45 9.10 ;
        RECT  3.15 5.55 7.25 6.05 ;
        RECT  6.20 2.55 6.90 3.25 ;
        RECT  6.20 9.75 6.90 10.45 ;
        RECT  6.55 5.55 7.25 6.25 ;
        RECT  6.20 2.75 8.25 3.25 ;
        RECT  7.55 6.65 8.05 10.25 ;
        RECT  7.75 2.75 8.05 10.25 ;
        RECT  6.20 9.75 8.05 10.25 ;
        RECT  7.75 2.75 8.25 7.15 ;
        RECT  9.05 4.25 9.80 4.95 ;
        RECT  9.20 6.45 9.90 7.15 ;
        RECT  7.55 6.65 9.90 7.15 ;
        RECT  9.05 4.45 10.90 4.95 ;
        RECT  10.40 4.45 10.90 8.35 ;
        RECT  10.05 7.65 10.90 8.35 ;
        RECT  12.05 6.45 12.75 7.15 ;
        RECT  10.40 6.65 12.75 7.15 ;
        RECT  13.25 2.75 13.75 8.35 ;
        RECT  12.75 7.65 13.75 8.35 ;
        RECT  13.25 5.50 15.35 6.00 ;
        RECT  14.10 2.55 14.80 3.25 ;
        RECT  13.25 2.75 14.80 3.25 ;
        RECT  14.65 5.50 15.35 6.20 ;
        RECT  15.65 4.25 16.35 4.95 ;
        RECT  15.85 4.25 16.35 10.50 ;
        RECT  15.60 7.65 16.35 10.50 ;
        RECT  15.60 9.80 16.65 10.50 ;
    END
END DLLRSX2
MACRO DLLRSX4
    CLASS CORE ;
    FOREIGN DLLRSX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  10.05 9.30 10.95 10.20 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  14.25 3.75 14.95 5.00 ;
        RECT  14.25 4.00 15.15 5.00 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  21.30 2.90 22.00 4.50 ;
        RECT  21.50 2.90 22.00 10.50 ;
        RECT  21.30 5.35 22.00 10.50 ;
        RECT  21.15 5.35 22.15 6.35 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  18.60 2.90 19.10 10.50 ;
        RECT  18.60 2.90 19.30 4.50 ;
        RECT  18.60 7.10 19.30 10.50 ;
        RECT  18.45 5.35 19.35 6.35 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.60 5.35 2.60 6.35 ;
        RECT  1.25 5.65 2.60 6.35 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.30 4.25 6.80 4.95 ;
        RECT  5.80 4.05 6.80 5.05 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.15 2.50 11.00 ;
        RECT  3.85 9.70 4.55 11.00 ;
        RECT  0.45 10.05 4.55 11.00 ;
        RECT  8.70 7.65 9.25 11.00 ;
        RECT  8.55 9.70 9.25 11.00 ;
        RECT  8.70 7.65 9.40 8.35 ;
        RECT  11.40 7.65 12.10 8.35 ;
        RECT  11.50 7.65 12.10 11.00 ;
        RECT  14.25 7.65 14.95 11.00 ;
        RECT  17.25 7.10 17.95 11.00 ;
        RECT  19.95 7.10 20.65 11.00 ;
        RECT  22.65 7.10 23.35 11.00 ;
        RECT  0.00 11.00 23.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.35 ;
        RECT  3.85 2.00 4.55 3.25 ;
        RECT  8.75 2.00 9.45 3.25 ;
        RECT  11.75 2.00 12.45 4.95 ;
        RECT  11.40 4.20 12.45 4.95 ;
        RECT  17.25 2.00 17.95 4.50 ;
        RECT  19.95 2.00 20.65 4.50 ;
        RECT  22.65 2.00 23.35 4.50 ;
        RECT  0.00 0.00 23.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.50 3.70 3.65 4.20 ;
        RECT  0.25 4.35 0.75 8.85 ;
        RECT  0.25 7.15 1.15 8.85 ;
        RECT  1.00 3.10 1.80 4.85 ;
        RECT  0.25 4.35 1.80 4.85 ;
        RECT  3.15 2.55 3.20 8.90 ;
        RECT  2.50 2.55 3.20 4.20 ;
        RECT  3.15 3.70 3.65 8.90 ;
        RECT  3.15 7.15 3.85 8.90 ;
        RECT  3.15 8.40 6.45 8.90 ;
        RECT  5.75 8.40 6.45 9.10 ;
        RECT  3.15 5.55 7.25 6.05 ;
        RECT  6.20 2.55 6.90 3.25 ;
        RECT  6.20 9.75 6.90 10.45 ;
        RECT  6.55 5.55 7.25 6.25 ;
        RECT  6.20 2.75 8.25 3.25 ;
        RECT  7.55 6.65 8.05 10.25 ;
        RECT  7.75 2.75 8.05 10.25 ;
        RECT  6.20 9.75 8.05 10.25 ;
        RECT  7.75 2.75 8.25 7.15 ;
        RECT  9.05 4.25 9.80 4.95 ;
        RECT  9.20 6.45 9.90 7.15 ;
        RECT  7.55 6.65 9.90 7.15 ;
        RECT  9.05 4.45 10.90 4.95 ;
        RECT  10.40 4.45 10.90 8.35 ;
        RECT  10.05 7.65 10.90 8.35 ;
        RECT  12.05 6.45 12.75 7.15 ;
        RECT  10.40 6.65 12.75 7.15 ;
        RECT  13.25 2.75 13.75 8.35 ;
        RECT  12.75 7.65 13.75 8.35 ;
        RECT  13.25 6.05 15.35 6.55 ;
        RECT  14.10 2.55 14.80 3.25 ;
        RECT  13.25 2.75 14.80 3.25 ;
        RECT  14.65 6.05 15.35 6.75 ;
        RECT  15.85 3.80 16.35 10.50 ;
        RECT  15.60 7.65 16.35 10.50 ;
        RECT  15.75 3.80 16.45 4.50 ;
        RECT  15.60 9.80 16.65 10.50 ;
    END
END DLLRSX4
MACRO DLLRX1
    CLASS CORE ;
    FOREIGN DLLRX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.35 15.15 6.35 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  17.15 3.75 17.95 4.45 ;
        RECT  17.05 5.35 17.95 6.35 ;
        RECT  17.35 3.75 17.95 8.90 ;
        RECT  17.15 7.15 17.95 8.90 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  19.85 3.75 20.35 8.90 ;
        RECT  19.85 3.75 20.55 4.45 ;
        RECT  19.85 7.15 20.55 8.90 ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.60 5.35 2.60 6.35 ;
        RECT  1.25 5.65 2.60 6.35 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.30 4.25 6.80 4.95 ;
        RECT  5.80 4.05 6.80 5.05 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.15 2.50 11.00 ;
        RECT  3.85 9.70 4.55 11.00 ;
        RECT  0.45 10.05 4.55 11.00 ;
        RECT  8.70 7.70 9.40 11.00 ;
        RECT  14.30 7.60 15.00 11.00 ;
        RECT  18.50 7.15 19.20 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.35 ;
        RECT  3.85 2.00 4.55 3.25 ;
        RECT  8.70 2.00 9.40 3.25 ;
        RECT  11.45 2.00 12.15 3.25 ;
        RECT  14.30 2.00 15.00 3.65 ;
        RECT  18.50 2.00 19.20 4.45 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.50 3.70 3.65 4.20 ;
        RECT  0.25 4.35 0.75 8.85 ;
        RECT  0.25 7.15 1.15 8.85 ;
        RECT  1.00 3.10 1.80 4.85 ;
        RECT  0.25 4.35 1.80 4.85 ;
        RECT  3.15 2.55 3.20 8.90 ;
        RECT  2.50 2.55 3.20 4.20 ;
        RECT  3.15 3.70 3.65 8.90 ;
        RECT  3.15 7.15 3.85 8.90 ;
        RECT  3.15 8.40 6.45 8.90 ;
        RECT  5.75 8.40 6.45 9.10 ;
        RECT  3.15 5.55 7.25 6.05 ;
        RECT  6.20 2.55 6.90 3.25 ;
        RECT  6.20 9.75 6.90 10.45 ;
        RECT  6.55 5.55 7.25 6.25 ;
        RECT  6.20 2.75 7.80 3.25 ;
        RECT  7.55 6.65 8.05 10.25 ;
        RECT  7.75 2.75 7.80 10.25 ;
        RECT  7.30 2.75 7.80 4.45 ;
        RECT  7.75 3.95 8.05 10.25 ;
        RECT  6.20 9.75 8.05 10.25 ;
        RECT  7.75 3.95 8.25 7.15 ;
        RECT  9.15 3.75 9.85 4.45 ;
        RECT  7.30 3.95 9.85 4.45 ;
        RECT  10.05 2.55 10.95 3.25 ;
        RECT  10.45 2.55 10.95 4.25 ;
        RECT  10.40 6.45 11.10 7.15 ;
        RECT  7.55 6.65 11.10 7.15 ;
        RECT  10.45 3.75 12.45 4.25 ;
        RECT  11.05 7.70 11.75 10.50 ;
        RECT  11.75 3.75 12.25 8.25 ;
        RECT  11.05 7.70 12.25 8.25 ;
        RECT  11.75 3.75 12.45 4.45 ;
        RECT  11.75 6.45 12.45 7.15 ;
        RECT  12.95 2.55 13.45 10.50 ;
        RECT  12.80 2.55 13.50 3.25 ;
        RECT  12.95 7.60 13.65 10.50 ;
        RECT  12.60 9.80 13.65 10.50 ;
        RECT  13.95 4.15 14.65 4.85 ;
        RECT  15.65 2.95 16.35 3.65 ;
        RECT  13.95 4.35 16.35 4.85 ;
        RECT  15.85 2.95 16.35 9.40 ;
        RECT  15.65 7.60 16.35 9.40 ;
    END
END DLLRX1
MACRO DLLRX2
    CLASS CORE ;
    FOREIGN DLLRX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.35 15.15 6.35 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  17.15 2.75 17.95 4.50 ;
        RECT  17.05 5.35 17.95 6.35 ;
        RECT  17.35 2.75 17.95 10.50 ;
        RECT  17.15 7.10 17.95 10.50 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  19.85 2.75 20.35 10.50 ;
        RECT  19.85 2.75 20.55 4.50 ;
        RECT  19.85 7.10 20.55 10.50 ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.60 5.35 2.60 6.35 ;
        RECT  1.25 5.65 2.60 6.35 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.30 4.25 6.80 4.95 ;
        RECT  5.80 4.05 6.80 5.05 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.15 2.50 11.00 ;
        RECT  3.85 9.70 4.55 11.00 ;
        RECT  0.45 10.05 4.55 11.00 ;
        RECT  8.70 7.70 9.40 11.00 ;
        RECT  14.30 7.60 15.00 11.00 ;
        RECT  18.50 7.10 19.20 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.35 ;
        RECT  3.85 2.00 4.55 3.25 ;
        RECT  8.70 2.00 9.40 3.25 ;
        RECT  11.45 2.00 12.15 3.25 ;
        RECT  14.30 2.00 15.00 3.65 ;
        RECT  18.50 2.00 19.20 4.50 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.50 3.70 3.65 4.20 ;
        RECT  0.25 4.35 0.75 8.85 ;
        RECT  0.25 7.15 1.15 8.85 ;
        RECT  1.00 3.10 1.80 4.85 ;
        RECT  0.25 4.35 1.80 4.85 ;
        RECT  3.15 2.55 3.20 8.90 ;
        RECT  2.50 2.55 3.20 4.20 ;
        RECT  3.15 3.70 3.65 8.90 ;
        RECT  3.15 7.15 3.85 8.90 ;
        RECT  3.15 8.40 6.45 8.90 ;
        RECT  5.75 8.40 6.45 9.10 ;
        RECT  3.15 5.55 7.25 6.05 ;
        RECT  6.20 2.55 6.90 3.25 ;
        RECT  6.20 9.75 6.90 10.45 ;
        RECT  6.55 5.55 7.25 6.25 ;
        RECT  6.20 2.75 7.80 3.25 ;
        RECT  7.55 6.65 8.05 10.25 ;
        RECT  7.75 2.75 7.80 10.25 ;
        RECT  7.30 2.75 7.80 4.45 ;
        RECT  7.75 3.95 8.05 10.25 ;
        RECT  6.20 9.75 8.05 10.25 ;
        RECT  7.75 3.95 8.25 7.15 ;
        RECT  9.15 3.75 9.85 4.45 ;
        RECT  7.30 3.95 9.85 4.45 ;
        RECT  10.05 2.55 10.95 3.25 ;
        RECT  10.45 2.55 10.95 4.25 ;
        RECT  10.40 6.45 11.10 7.15 ;
        RECT  7.55 6.65 11.10 7.15 ;
        RECT  10.45 3.75 12.45 4.25 ;
        RECT  11.05 7.70 11.75 10.50 ;
        RECT  11.75 3.75 12.25 8.25 ;
        RECT  11.05 7.70 12.25 8.25 ;
        RECT  11.75 3.75 12.45 4.45 ;
        RECT  11.75 6.45 12.45 7.15 ;
        RECT  12.95 2.55 13.45 10.50 ;
        RECT  12.80 2.55 13.50 3.25 ;
        RECT  12.95 7.60 13.65 10.50 ;
        RECT  12.60 9.80 13.65 10.50 ;
        RECT  13.95 4.15 14.65 4.85 ;
        RECT  15.65 2.95 16.35 3.65 ;
        RECT  13.95 4.35 16.35 4.85 ;
        RECT  15.85 2.95 16.35 9.40 ;
        RECT  15.65 7.60 16.35 9.40 ;
    END
END DLLRX2
MACRO DLLRX4
    CLASS CORE ;
    FOREIGN DLLRX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.35 15.15 6.35 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  18.60 2.90 19.10 10.50 ;
        RECT  18.60 2.90 19.30 4.50 ;
        RECT  18.60 7.10 19.30 10.50 ;
        RECT  18.45 5.35 19.35 6.35 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  21.30 2.90 22.00 4.50 ;
        RECT  21.50 2.90 22.00 10.50 ;
        RECT  21.30 5.35 22.00 10.50 ;
        RECT  21.25 5.35 22.15 6.35 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.60 5.35 2.60 6.35 ;
        RECT  1.25 5.65 2.60 6.35 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.30 4.25 6.80 4.95 ;
        RECT  5.80 4.05 6.80 5.05 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.15 2.50 11.00 ;
        RECT  3.85 9.70 4.55 11.00 ;
        RECT  0.45 10.05 4.55 11.00 ;
        RECT  8.70 7.70 9.40 11.00 ;
        RECT  14.30 7.60 15.00 11.00 ;
        RECT  17.25 7.10 17.95 11.00 ;
        RECT  19.95 7.10 20.65 11.00 ;
        RECT  22.65 7.10 23.35 11.00 ;
        RECT  0.00 11.00 23.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.35 ;
        RECT  3.85 2.00 4.55 3.25 ;
        RECT  8.70 2.00 9.40 3.25 ;
        RECT  11.45 2.00 12.15 3.25 ;
        RECT  14.30 2.00 15.00 3.65 ;
        RECT  17.25 2.00 17.95 4.50 ;
        RECT  19.95 2.00 20.65 4.50 ;
        RECT  22.65 2.00 23.35 4.50 ;
        RECT  0.00 0.00 23.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.50 3.70 3.65 4.20 ;
        RECT  0.25 4.35 0.75 8.85 ;
        RECT  0.25 7.15 1.15 8.85 ;
        RECT  1.00 3.10 1.80 4.85 ;
        RECT  0.25 4.35 1.80 4.85 ;
        RECT  3.15 2.55 3.20 8.90 ;
        RECT  2.50 2.55 3.20 4.20 ;
        RECT  3.15 3.70 3.65 8.90 ;
        RECT  3.15 7.15 3.85 8.90 ;
        RECT  3.15 8.40 6.45 8.90 ;
        RECT  5.75 8.40 6.45 9.10 ;
        RECT  3.15 5.55 7.25 6.05 ;
        RECT  6.20 2.55 6.90 3.25 ;
        RECT  6.20 9.75 6.90 10.45 ;
        RECT  6.55 5.55 7.25 6.25 ;
        RECT  6.20 2.75 7.80 3.25 ;
        RECT  7.55 6.65 8.05 10.25 ;
        RECT  7.75 2.75 7.80 10.25 ;
        RECT  7.30 2.75 7.80 4.45 ;
        RECT  7.75 3.95 8.05 10.25 ;
        RECT  6.20 9.75 8.05 10.25 ;
        RECT  7.75 3.95 8.25 7.15 ;
        RECT  9.15 3.75 9.85 4.45 ;
        RECT  7.30 3.95 9.85 4.45 ;
        RECT  10.05 2.55 10.95 3.25 ;
        RECT  10.45 2.55 10.95 4.25 ;
        RECT  10.40 6.45 11.10 7.15 ;
        RECT  7.55 6.65 11.10 7.15 ;
        RECT  10.45 3.75 12.45 4.25 ;
        RECT  11.05 7.70 11.75 10.50 ;
        RECT  11.75 3.75 12.25 8.25 ;
        RECT  11.05 7.70 12.25 8.25 ;
        RECT  11.75 3.75 12.45 4.45 ;
        RECT  11.75 6.45 12.45 7.15 ;
        RECT  12.95 2.55 13.45 10.50 ;
        RECT  12.80 2.55 13.50 3.25 ;
        RECT  12.95 7.60 13.65 10.50 ;
        RECT  12.60 9.80 13.65 10.50 ;
        RECT  13.95 4.15 14.65 4.85 ;
        RECT  15.65 2.95 16.35 3.65 ;
        RECT  13.95 4.35 16.35 4.85 ;
        RECT  15.85 2.95 16.35 9.40 ;
        RECT  15.65 7.60 16.35 9.40 ;
    END
END DLLRX4
MACRO DLLSX1
    CLASS CORE ;
    FOREIGN DLLSX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  11.15 4.25 12.35 4.95 ;
        RECT  11.45 4.10 12.35 5.00 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  17.05 3.75 17.60 9.65 ;
        RECT  17.05 3.75 17.75 4.45 ;
        RECT  17.05 7.90 17.75 9.65 ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  14.35 3.75 15.15 4.45 ;
        RECT  14.25 5.40 15.15 6.30 ;
        RECT  14.65 3.75 15.15 9.65 ;
        RECT  14.35 8.00 15.15 9.65 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.15 8.25 ;
        RECT  1.45 7.55 2.15 8.25 ;
        RECT  1.65 6.70 2.55 7.60 ;
        RECT  1.45 7.55 2.55 7.60 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 8.00 5.35 8.90 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.75 2.50 11.00 ;
        RECT  4.80 9.40 5.50 11.00 ;
        RECT  8.80 7.35 9.50 8.05 ;
        RECT  9.00 7.35 9.50 9.05 ;
        RECT  9.50 8.55 10.20 11.00 ;
        RECT  11.50 7.35 12.00 9.05 ;
        RECT  9.00 8.55 12.00 9.05 ;
        RECT  11.50 7.35 12.20 8.05 ;
        RECT  15.70 7.90 16.40 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.60 ;
        RECT  1.80 4.00 3.50 4.60 ;
        RECT  2.80 4.00 3.50 5.85 ;
        RECT  7.65 2.00 8.35 4.05 ;
        RECT  11.50 2.00 12.20 3.60 ;
        RECT  15.70 2.00 16.40 4.45 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  12.85 3.15 13.75 3.65 ;
        RECT  0.25 8.75 1.15 9.25 ;
        RECT  0.45 2.55 0.75 10.45 ;
        RECT  0.25 2.55 0.75 9.25 ;
        RECT  0.25 2.55 1.15 3.25 ;
        RECT  0.45 8.75 1.15 10.45 ;
        RECT  0.25 5.45 2.30 6.15 ;
        RECT  3.15 6.75 3.65 10.45 ;
        RECT  3.15 2.55 3.85 3.25 ;
        RECT  3.15 8.75 3.85 10.45 ;
        RECT  3.15 2.75 4.50 3.25 ;
        RECT  4.00 2.75 4.50 7.25 ;
        RECT  5.30 3.45 6.00 5.85 ;
        RECT  5.15 5.10 6.00 5.85 ;
        RECT  3.15 6.75 6.90 7.25 ;
        RECT  6.20 6.75 6.90 7.45 ;
        RECT  5.15 5.35 7.90 5.85 ;
        RECT  7.40 5.35 7.90 10.45 ;
        RECT  7.15 9.75 7.90 10.45 ;
        RECT  7.40 6.15 9.65 6.85 ;
        RECT  9.15 2.95 9.85 3.65 ;
        RECT  9.15 3.15 10.65 3.65 ;
        RECT  10.15 3.15 10.65 8.05 ;
        RECT  10.15 5.75 10.85 8.05 ;
        RECT  10.85 9.75 11.55 10.45 ;
        RECT  11.95 5.55 12.65 6.25 ;
        RECT  10.15 5.75 12.65 6.25 ;
        RECT  13.25 2.95 13.55 10.25 ;
        RECT  12.85 2.95 13.55 3.65 ;
        RECT  13.25 3.15 13.75 10.25 ;
        RECT  10.85 9.75 13.75 10.25 ;
        RECT  13.25 6.80 14.15 7.50 ;
    END
END DLLSX1
MACRO DLLSX2
    CLASS CORE ;
    FOREIGN DLLSX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  11.15 4.25 12.35 4.95 ;
        RECT  11.45 4.10 12.35 5.00 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  17.05 2.70 17.60 10.50 ;
        RECT  17.05 2.70 17.75 4.50 ;
        RECT  17.05 7.10 17.75 10.50 ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  14.35 2.70 15.15 4.50 ;
        RECT  14.25 5.40 15.15 6.30 ;
        RECT  14.65 2.70 15.15 10.50 ;
        RECT  14.35 7.10 15.15 10.50 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.15 8.25 ;
        RECT  1.45 7.55 2.15 8.25 ;
        RECT  1.65 6.70 2.55 7.60 ;
        RECT  1.45 7.55 2.55 7.60 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 8.00 5.35 8.90 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.75 2.50 11.00 ;
        RECT  4.80 9.40 5.50 11.00 ;
        RECT  8.45 7.35 9.15 8.05 ;
        RECT  8.60 7.35 9.15 9.05 ;
        RECT  9.50 8.55 10.20 11.00 ;
        RECT  11.15 7.35 11.65 9.05 ;
        RECT  8.60 8.55 11.65 9.05 ;
        RECT  11.15 7.35 11.85 8.05 ;
        RECT  15.70 7.10 16.40 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.60 ;
        RECT  1.80 4.00 3.50 4.60 ;
        RECT  2.80 4.00 3.50 5.85 ;
        RECT  7.65 2.00 8.35 4.05 ;
        RECT  11.50 2.00 12.20 3.50 ;
        RECT  15.70 2.00 16.40 4.50 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  9.15 3.05 10.30 3.55 ;
        RECT  12.85 3.05 13.75 3.55 ;
        RECT  0.25 8.75 1.15 9.25 ;
        RECT  0.45 2.55 0.75 10.45 ;
        RECT  0.25 2.55 0.75 9.25 ;
        RECT  0.25 2.55 1.15 3.25 ;
        RECT  0.45 8.75 1.15 10.45 ;
        RECT  0.25 5.45 2.30 6.15 ;
        RECT  3.15 6.75 3.65 10.45 ;
        RECT  3.15 2.55 3.85 3.25 ;
        RECT  3.15 8.75 3.85 10.45 ;
        RECT  3.15 2.75 4.50 3.25 ;
        RECT  4.00 2.75 4.50 7.25 ;
        RECT  5.30 3.45 6.00 5.85 ;
        RECT  5.15 5.10 6.00 5.85 ;
        RECT  3.15 6.75 6.90 7.25 ;
        RECT  6.20 6.75 6.90 7.45 ;
        RECT  5.15 5.35 7.90 5.85 ;
        RECT  7.40 5.35 7.90 10.45 ;
        RECT  7.15 9.75 7.90 10.45 ;
        RECT  7.40 6.15 9.30 6.85 ;
        RECT  9.80 2.85 9.85 8.05 ;
        RECT  9.15 2.85 9.85 3.55 ;
        RECT  9.80 3.05 10.30 8.05 ;
        RECT  9.80 5.70 10.50 8.05 ;
        RECT  10.85 9.75 11.55 10.45 ;
        RECT  11.95 5.50 12.65 6.20 ;
        RECT  9.80 5.70 12.65 6.20 ;
        RECT  13.25 2.85 13.55 10.25 ;
        RECT  12.85 2.85 13.55 3.55 ;
        RECT  13.25 3.05 13.75 10.25 ;
        RECT  10.85 9.75 13.75 10.25 ;
        RECT  13.15 6.55 13.85 7.25 ;
    END
END DLLSX2
MACRO DLLSX4
    CLASS CORE ;
    FOREIGN DLLSX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  11.15 4.25 12.35 4.95 ;
        RECT  11.45 4.10 12.35 5.00 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  18.50 2.90 19.20 4.50 ;
        RECT  18.70 2.90 19.20 10.50 ;
        RECT  18.50 5.35 19.20 10.50 ;
        RECT  18.35 5.35 19.35 6.35 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  15.80 2.90 16.30 10.50 ;
        RECT  15.80 2.90 16.50 4.50 ;
        RECT  15.80 7.10 16.50 10.50 ;
        RECT  15.65 5.35 16.55 6.35 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.15 8.25 ;
        RECT  1.45 7.55 2.15 8.25 ;
        RECT  1.65 6.70 2.55 7.60 ;
        RECT  1.45 7.55 2.55 7.60 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 8.00 5.35 8.90 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.75 2.50 11.00 ;
        RECT  4.80 9.40 5.50 11.00 ;
        RECT  8.45 7.35 9.15 8.05 ;
        RECT  8.60 7.35 9.15 9.05 ;
        RECT  9.50 8.55 10.20 11.00 ;
        RECT  11.15 7.35 11.65 9.05 ;
        RECT  8.60 8.55 11.65 9.05 ;
        RECT  11.15 7.35 11.85 8.05 ;
        RECT  14.45 7.10 15.15 11.00 ;
        RECT  17.15 7.10 17.85 11.00 ;
        RECT  19.85 7.10 20.55 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.60 ;
        RECT  1.80 4.00 3.50 4.60 ;
        RECT  2.80 4.00 3.50 5.85 ;
        RECT  7.65 2.00 8.35 4.05 ;
        RECT  11.50 2.00 12.20 3.50 ;
        RECT  14.45 2.00 15.15 4.50 ;
        RECT  17.15 2.00 17.85 4.50 ;
        RECT  19.85 2.00 20.55 4.50 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  9.15 3.05 10.30 3.55 ;
        RECT  12.85 3.05 13.75 3.55 ;
        RECT  0.25 8.75 1.15 9.25 ;
        RECT  0.45 2.55 0.75 10.45 ;
        RECT  0.25 2.55 0.75 9.25 ;
        RECT  0.25 2.55 1.15 3.25 ;
        RECT  0.45 8.75 1.15 10.45 ;
        RECT  0.25 5.45 2.30 6.15 ;
        RECT  3.15 6.75 3.65 10.45 ;
        RECT  3.15 2.55 3.85 3.25 ;
        RECT  3.15 8.75 3.85 10.45 ;
        RECT  3.15 2.75 4.50 3.25 ;
        RECT  4.00 2.75 4.50 7.25 ;
        RECT  5.30 3.45 6.00 5.85 ;
        RECT  5.15 5.10 6.00 5.85 ;
        RECT  3.15 6.75 6.90 7.25 ;
        RECT  6.20 6.75 6.90 7.45 ;
        RECT  5.15 5.35 7.90 5.85 ;
        RECT  7.40 5.35 7.90 10.45 ;
        RECT  7.15 9.75 7.90 10.45 ;
        RECT  7.40 6.15 9.30 6.85 ;
        RECT  9.80 2.85 9.85 8.05 ;
        RECT  9.15 2.85 9.85 3.55 ;
        RECT  9.80 3.05 10.30 8.05 ;
        RECT  9.80 5.70 10.50 8.05 ;
        RECT  10.85 9.75 11.55 10.45 ;
        RECT  11.95 5.50 12.65 6.20 ;
        RECT  9.80 5.70 12.65 6.20 ;
        RECT  13.25 2.85 13.55 10.25 ;
        RECT  12.85 2.85 13.55 3.55 ;
        RECT  13.25 3.05 13.75 10.25 ;
        RECT  10.85 9.75 13.75 10.25 ;
        RECT  13.15 6.55 13.85 7.25 ;
    END
END DLLSX4
MACRO DLLX1
    CLASS CORE ;
    FOREIGN DLLX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  14.25 3.55 14.80 8.90 ;
        RECT  14.25 3.55 14.95 4.25 ;
        RECT  14.25 7.15 14.95 8.90 ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.55 3.55 12.35 4.25 ;
        RECT  11.45 5.40 12.35 6.30 ;
        RECT  11.85 3.55 12.35 8.90 ;
        RECT  11.55 7.25 12.35 8.90 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.15 8.25 ;
        RECT  1.45 7.55 2.15 8.25 ;
        RECT  1.65 6.70 2.55 7.60 ;
        RECT  1.45 7.55 2.55 7.60 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 8.00 5.35 8.90 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.75 2.50 11.00 ;
        RECT  4.80 9.40 5.50 11.00 ;
        RECT  8.45 6.90 9.15 11.00 ;
        RECT  8.45 10.30 10.40 11.00 ;
        RECT  12.90 7.15 13.60 11.00 ;
        RECT  11.35 10.10 14.95 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.60 ;
        RECT  1.80 4.00 3.50 4.60 ;
        RECT  2.80 4.00 3.50 5.85 ;
        RECT  7.65 2.00 8.35 4.20 ;
        RECT  12.90 2.00 13.60 4.25 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 2.55 0.95 10.45 ;
        RECT  0.45 2.55 1.15 3.25 ;
        RECT  0.45 8.75 1.15 10.45 ;
        RECT  0.45 5.45 2.30 6.15 ;
        RECT  3.15 6.75 3.65 10.45 ;
        RECT  3.15 2.55 3.85 3.25 ;
        RECT  3.15 8.75 3.85 10.45 ;
        RECT  3.15 2.75 4.50 3.25 ;
        RECT  4.00 2.75 4.50 7.25 ;
        RECT  5.30 3.60 5.85 5.85 ;
        RECT  5.15 5.10 5.85 5.85 ;
        RECT  5.30 3.60 6.00 4.30 ;
        RECT  3.15 6.75 6.90 7.25 ;
        RECT  6.20 6.75 6.90 7.45 ;
        RECT  7.40 5.35 7.90 10.50 ;
        RECT  7.15 9.80 7.90 10.50 ;
        RECT  5.15 5.35 9.25 5.85 ;
        RECT  8.55 5.35 9.25 6.05 ;
        RECT  9.00 3.60 10.50 4.30 ;
        RECT  10.00 2.50 10.50 9.75 ;
        RECT  9.80 6.90 10.50 9.75 ;
        RECT  10.00 2.50 10.75 3.20 ;
        RECT  9.80 9.05 10.85 9.75 ;
    END
END DLLX1
MACRO DLLX2
    CLASS CORE ;
    FOREIGN DLLX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  14.25 2.75 14.80 10.50 ;
        RECT  14.25 2.75 14.95 4.50 ;
        RECT  14.25 7.10 14.95 10.50 ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.55 2.70 12.35 4.30 ;
        RECT  11.45 5.40 12.35 6.30 ;
        RECT  11.85 2.70 12.35 10.50 ;
        RECT  11.55 7.10 12.35 10.50 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.15 8.25 ;
        RECT  1.45 7.55 2.15 8.25 ;
        RECT  1.65 6.70 2.55 7.60 ;
        RECT  1.45 7.55 2.55 7.60 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 8.00 5.35 8.90 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.75 2.50 11.00 ;
        RECT  4.80 9.40 5.50 11.00 ;
        RECT  8.45 6.90 9.15 11.00 ;
        RECT  8.45 10.30 10.40 11.00 ;
        RECT  12.90 7.10 13.60 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.60 ;
        RECT  1.80 4.00 3.50 4.60 ;
        RECT  2.80 4.00 3.50 5.85 ;
        RECT  7.65 2.00 8.35 4.20 ;
        RECT  12.90 2.00 13.60 4.50 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 2.55 0.95 10.45 ;
        RECT  0.45 2.55 1.15 3.25 ;
        RECT  0.45 8.75 1.15 10.45 ;
        RECT  0.45 5.45 2.30 6.15 ;
        RECT  3.15 6.75 3.65 10.45 ;
        RECT  3.15 2.55 3.85 3.25 ;
        RECT  3.15 8.75 3.85 10.45 ;
        RECT  3.15 2.75 4.50 3.25 ;
        RECT  4.00 2.75 4.50 7.25 ;
        RECT  5.30 3.60 5.85 5.85 ;
        RECT  5.15 5.10 5.85 5.85 ;
        RECT  5.30 3.60 6.00 4.30 ;
        RECT  3.15 6.75 6.90 7.25 ;
        RECT  6.20 6.75 6.90 7.45 ;
        RECT  7.40 5.35 7.90 10.50 ;
        RECT  7.15 9.80 7.90 10.50 ;
        RECT  5.15 5.35 9.25 5.85 ;
        RECT  8.55 5.35 9.25 6.05 ;
        RECT  9.00 3.60 10.50 4.30 ;
        RECT  10.00 2.50 10.50 9.75 ;
        RECT  9.80 7.10 10.50 9.75 ;
        RECT  10.00 2.50 10.75 3.20 ;
        RECT  9.80 9.05 10.85 9.75 ;
    END
END DLLX2
MACRO DLLX4
    CLASS CORE ;
    FOREIGN DLLX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  15.70 2.90 16.40 4.50 ;
        RECT  15.90 2.90 16.40 10.50 ;
        RECT  15.70 5.35 16.40 10.50 ;
        RECT  15.55 5.35 16.55 6.35 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  13.00 2.90 13.50 10.50 ;
        RECT  13.00 2.90 13.70 4.50 ;
        RECT  13.00 7.10 13.70 10.50 ;
        RECT  12.85 5.35 13.75 6.35 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.15 8.25 ;
        RECT  1.45 7.55 2.15 8.25 ;
        RECT  1.65 6.70 2.55 7.60 ;
        RECT  1.45 7.55 2.55 7.60 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 8.00 5.35 8.90 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.75 2.50 11.00 ;
        RECT  4.80 9.40 5.50 11.00 ;
        RECT  8.45 6.90 9.15 11.00 ;
        RECT  8.45 10.30 10.40 11.00 ;
        RECT  11.65 7.10 12.35 11.00 ;
        RECT  14.35 7.10 15.05 11.00 ;
        RECT  17.05 7.10 17.75 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.60 ;
        RECT  1.80 4.00 3.50 4.60 ;
        RECT  2.80 4.00 3.50 5.85 ;
        RECT  7.65 2.00 8.35 4.20 ;
        RECT  11.65 2.00 12.35 4.30 ;
        RECT  14.35 2.00 15.05 4.50 ;
        RECT  17.05 2.00 17.75 4.50 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 2.55 0.95 10.45 ;
        RECT  0.45 2.55 1.15 3.25 ;
        RECT  0.45 8.75 1.15 10.45 ;
        RECT  0.45 5.45 2.30 6.15 ;
        RECT  3.15 6.75 3.65 10.45 ;
        RECT  3.15 2.55 3.85 3.25 ;
        RECT  3.15 8.75 3.85 10.45 ;
        RECT  3.15 2.75 4.50 3.25 ;
        RECT  4.00 2.75 4.50 7.25 ;
        RECT  5.30 3.60 5.85 5.85 ;
        RECT  5.15 5.10 5.85 5.85 ;
        RECT  5.30 3.60 6.00 4.30 ;
        RECT  3.15 6.75 6.90 7.25 ;
        RECT  6.20 6.75 6.90 7.45 ;
        RECT  7.40 5.35 7.90 10.50 ;
        RECT  7.15 9.80 7.90 10.50 ;
        RECT  5.15 5.35 9.25 5.85 ;
        RECT  8.55 5.35 9.25 6.05 ;
        RECT  9.00 3.60 10.50 4.30 ;
        RECT  10.00 2.50 10.50 9.75 ;
        RECT  9.80 7.10 10.50 9.75 ;
        RECT  10.00 2.50 10.75 3.20 ;
        RECT  9.80 9.05 10.85 9.75 ;
    END
END DLLX4
MACRO DLY1X1
    CLASS CORE ;
    FOREIGN DLY1X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.65 2.85 9.35 5.00 ;
        RECT  8.85 2.85 9.35 8.90 ;
        RECT  8.65 7.05 9.35 8.90 ;
        RECT  8.65 4.10 9.55 5.00 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.05 2.50 11.00 ;
        RECT  7.30 7.95 8.00 11.00 ;
        RECT  0.45 10.30 9.35 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.55 2.00 7.85 2.90 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.75 1.15 4.45 ;
        RECT  0.45 7.10 1.15 8.90 ;
        RECT  0.45 3.90 3.30 4.45 ;
        RECT  2.80 3.90 3.30 7.60 ;
        RECT  0.45 7.10 3.30 7.60 ;
        RECT  2.80 4.75 3.50 6.65 ;
        RECT  3.80 3.70 4.60 4.40 ;
        RECT  4.10 3.70 4.60 7.85 ;
        RECT  3.90 7.10 4.60 7.85 ;
        RECT  5.40 7.00 5.90 9.30 ;
        RECT  5.20 8.55 5.90 9.30 ;
        RECT  5.30 3.75 6.00 4.45 ;
        RECT  6.30 4.90 7.00 6.50 ;
        RECT  4.10 6.00 7.00 6.50 ;
        RECT  5.30 3.95 8.15 4.45 ;
        RECT  7.65 3.95 8.15 7.50 ;
        RECT  5.40 7.00 8.15 7.50 ;
        RECT  7.65 5.60 8.40 6.30 ;
    END
END DLY1X1
MACRO DLY2X1
    CLASS CORE ;
    FOREIGN DLY2X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  14.35 2.85 14.90 8.90 ;
        RECT  14.20 7.10 14.90 8.90 ;
        RECT  14.25 2.85 14.95 5.00 ;
        RECT  14.25 4.10 15.15 5.00 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.05 2.50 11.00 ;
        RECT  7.40 7.90 8.10 11.00 ;
        RECT  12.85 7.95 13.55 11.00 ;
        RECT  0.45 10.15 14.95 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.55 2.00 4.20 2.90 ;
        RECT  7.35 2.00 8.05 3.35 ;
        RECT  11.05 2.00 13.45 2.90 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.75 1.15 4.45 ;
        RECT  0.45 7.10 1.15 8.90 ;
        RECT  0.45 3.95 3.30 4.45 ;
        RECT  2.80 3.95 3.30 7.60 ;
        RECT  0.45 7.10 3.30 7.60 ;
        RECT  2.80 4.85 3.50 6.65 ;
        RECT  3.80 3.75 4.60 4.45 ;
        RECT  4.10 3.75 4.60 9.30 ;
        RECT  3.90 8.60 4.60 9.30 ;
        RECT  5.30 3.75 6.00 4.45 ;
        RECT  5.30 6.95 6.00 7.95 ;
        RECT  4.10 4.90 6.95 5.40 ;
        RECT  6.25 4.90 6.95 6.50 ;
        RECT  5.30 3.95 8.90 4.45 ;
        RECT  8.40 3.95 8.90 7.45 ;
        RECT  5.30 6.95 8.90 7.45 ;
        RECT  8.40 4.85 9.10 6.60 ;
        RECT  9.40 3.75 10.20 4.45 ;
        RECT  9.70 3.75 10.20 7.90 ;
        RECT  9.50 7.20 10.20 7.90 ;
        RECT  10.95 7.00 11.45 9.30 ;
        RECT  10.75 8.60 11.45 9.30 ;
        RECT  10.90 3.75 11.60 4.45 ;
        RECT  11.90 4.90 12.60 6.55 ;
        RECT  9.70 6.05 12.60 6.55 ;
        RECT  10.90 3.95 13.70 4.45 ;
        RECT  13.20 3.95 13.70 7.50 ;
        RECT  10.95 7.00 13.70 7.50 ;
        RECT  13.20 5.70 13.90 6.40 ;
    END
END DLY2X1
MACRO DLY4X1
    CLASS CORE ;
    FOREIGN DLY4X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  15.65 2.85 16.35 5.00 ;
        RECT  15.85 2.85 16.35 8.90 ;
        RECT  15.65 7.10 16.35 8.90 ;
        RECT  15.65 4.10 16.55 5.00 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.05 2.50 11.00 ;
        RECT  14.30 8.15 15.00 11.00 ;
        RECT  0.45 10.30 16.35 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.55 2.00 8.25 2.90 ;
        RECT  10.55 2.00 13.35 3.35 ;
        RECT  14.15 2.00 14.85 3.40 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.75 1.15 4.45 ;
        RECT  0.45 7.10 1.15 8.90 ;
        RECT  0.45 3.95 2.15 4.45 ;
        RECT  1.65 3.95 2.15 7.60 ;
        RECT  0.45 7.10 2.15 7.60 ;
        RECT  1.65 5.65 7.10 6.35 ;
        RECT  7.45 3.80 8.15 4.50 ;
        RECT  7.60 3.80 8.10 7.80 ;
        RECT  7.40 7.10 8.10 7.80 ;
        RECT  7.60 3.80 8.15 6.55 ;
        RECT  8.90 7.00 9.40 9.15 ;
        RECT  8.70 8.45 9.40 9.15 ;
        RECT  9.05 2.70 9.75 4.50 ;
        RECT  9.70 5.80 14.10 6.55 ;
        RECT  7.60 6.05 14.10 6.55 ;
        RECT  9.05 4.00 15.10 4.50 ;
        RECT  14.60 4.00 15.10 7.50 ;
        RECT  8.90 7.00 15.10 7.50 ;
        RECT  14.60 5.40 15.40 6.10 ;
    END
END DLY4X1
MACRO DLY8X1
    CLASS CORE ;
    FOREIGN DLY8X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 29.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  28.25 2.85 28.95 5.00 ;
        RECT  28.45 2.85 28.95 8.90 ;
        RECT  28.25 7.10 28.95 8.90 ;
        RECT  28.25 4.10 29.15 5.00 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.05 2.50 11.00 ;
        RECT  14.30 7.95 15.00 11.00 ;
        RECT  26.90 7.95 27.60 11.00 ;
        RECT  0.45 10.70 28.95 11.00 ;
        RECT  0.00 11.00 29.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.55 2.00 27.45 2.90 ;
        RECT  0.00 0.00 29.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.75 1.15 4.45 ;
        RECT  0.45 7.10 1.15 8.90 ;
        RECT  0.45 3.95 2.10 4.45 ;
        RECT  1.60 3.95 2.10 7.60 ;
        RECT  0.45 7.10 2.10 7.60 ;
        RECT  1.60 5.65 7.10 6.35 ;
        RECT  7.30 3.75 8.15 4.45 ;
        RECT  7.60 3.75 8.10 7.80 ;
        RECT  7.40 7.10 8.10 7.80 ;
        RECT  7.60 3.75 8.15 6.40 ;
        RECT  8.90 7.00 9.40 9.15 ;
        RECT  8.70 8.45 9.40 9.15 ;
        RECT  8.80 3.75 9.50 4.45 ;
        RECT  9.70 5.70 14.10 6.40 ;
        RECT  7.60 5.90 14.10 6.40 ;
        RECT  8.80 3.95 15.70 4.45 ;
        RECT  15.20 3.95 15.70 7.50 ;
        RECT  8.90 7.00 15.70 7.50 ;
        RECT  15.20 5.65 19.60 6.35 ;
        RECT  19.90 3.75 20.60 4.45 ;
        RECT  20.10 3.75 20.60 7.80 ;
        RECT  19.90 7.10 20.60 7.80 ;
        RECT  21.50 7.00 22.00 9.10 ;
        RECT  21.30 8.40 22.00 9.10 ;
        RECT  21.40 3.75 22.10 4.45 ;
        RECT  22.30 5.70 26.70 6.40 ;
        RECT  20.10 5.90 26.70 6.40 ;
        RECT  21.40 3.95 27.70 4.45 ;
        RECT  27.20 3.95 27.70 7.50 ;
        RECT  21.50 7.00 27.70 7.50 ;
        RECT  27.20 5.40 28.00 6.10 ;
    END
END DLY8X1
MACRO EN2X1
    CLASS CORE ;
    FOREIGN EN2X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  2.05 4.40 2.55 7.10 ;
        RECT  3.15 2.50 3.85 4.90 ;
        RECT  2.05 4.40 3.85 4.90 ;
        RECT  2.05 6.60 5.40 7.10 ;
        RECT  4.90 6.60 5.40 10.50 ;
        RECT  4.90 7.50 5.60 10.50 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.80 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.75 6.10 ;
        RECT  3.05 5.40 6.75 5.90 ;
        RECT  5.45 5.40 6.75 6.10 ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.80 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.40 7.60 4.10 11.00 ;
        RECT  7.25 7.50 7.95 11.00 ;
        RECT  0.00 11.00 8.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  5.90 2.00 6.60 3.90 ;
        RECT  0.00 0.00 8.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.65 3.40 1.15 8.05 ;
        RECT  0.65 7.55 2.60 8.05 ;
        RECT  1.90 7.55 2.60 8.30 ;
        RECT  1.40 3.20 2.10 3.90 ;
        RECT  0.65 3.40 2.10 3.90 ;
        RECT  2.10 7.55 2.60 10.00 ;
        RECT  1.10 9.30 2.90 10.00 ;
        RECT  4.50 2.50 5.20 4.10 ;
        RECT  4.70 2.50 5.20 4.90 ;
        RECT  7.25 2.50 7.75 4.90 ;
        RECT  4.70 4.40 7.75 4.90 ;
        RECT  7.25 2.50 7.95 4.10 ;
    END
END EN2X1
MACRO EN2X2
    CLASS CORE ;
    FOREIGN EN2X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.30 6.50 4.80 10.55 ;
        RECT  4.10 7.55 4.80 10.55 ;
        RECT  5.95 3.40 6.65 7.00 ;
        RECT  5.85 5.40 6.75 7.00 ;
        RECT  4.30 6.50 7.80 7.00 ;
        RECT  7.10 6.50 7.80 9.60 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.40 9.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.75 7.60 3.45 11.00 ;
        RECT  9.95 7.70 10.65 11.00 ;
        RECT  12.65 7.15 13.35 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.90 2.00 3.60 4.45 ;
        RECT  8.80 2.00 9.50 4.00 ;
        RECT  11.50 2.00 12.20 4.00 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.55 3.75 1.25 4.45 ;
        RECT  0.70 3.75 1.25 6.00 ;
        RECT  1.25 7.45 1.95 8.15 ;
        RECT  1.40 5.50 1.95 10.55 ;
        RECT  1.25 9.85 1.95 10.55 ;
        RECT  0.70 5.50 4.35 6.00 ;
        RECT  3.65 5.35 4.35 6.05 ;
        RECT  4.60 2.45 5.30 4.80 ;
        RECT  5.75 7.60 6.45 10.55 ;
        RECT  4.60 2.45 8.15 2.95 ;
        RECT  7.45 2.45 8.15 4.95 ;
        RECT  8.45 6.75 9.15 10.55 ;
        RECT  5.75 10.05 9.15 10.55 ;
        RECT  10.15 2.45 10.85 4.95 ;
        RECT  8.45 6.75 12.00 7.25 ;
        RECT  11.30 6.75 12.00 10.55 ;
        RECT  12.85 2.45 13.35 4.95 ;
        RECT  7.45 4.45 13.35 4.95 ;
        RECT  12.85 2.45 13.55 4.05 ;
    END
END EN2X2
MACRO EN2X3
    CLASS CORE ;
    FOREIGN EN2X3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  3.40 2.55 4.10 5.10 ;
        RECT  4.75 6.75 5.45 10.05 ;
        RECT  3.75 8.10 5.45 10.05 ;
        RECT  3.40 4.60 6.80 5.10 ;
        RECT  6.10 3.40 6.80 7.25 ;
        RECT  5.85 4.60 6.80 7.25 ;
        RECT  4.75 6.75 8.15 7.25 ;
        RECT  7.45 6.75 8.15 9.60 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 7.00 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 7.00 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.40 7.10 3.10 11.00 ;
        RECT  2.40 10.70 4.30 11.00 ;
        RECT  10.15 7.70 10.85 11.00 ;
        RECT  12.85 7.15 13.55 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  8.80 2.00 9.50 4.00 ;
        RECT  11.50 2.00 12.20 4.00 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.90 3.60 1.40 10.55 ;
        RECT  0.90 7.45 1.60 8.15 ;
        RECT  0.90 9.85 1.60 10.55 ;
        RECT  0.90 3.60 1.65 4.30 ;
        RECT  0.90 5.55 4.55 6.05 ;
        RECT  3.85 5.55 4.55 6.25 ;
        RECT  4.75 2.45 5.45 4.15 ;
        RECT  6.10 7.70 6.80 10.55 ;
        RECT  4.75 2.45 8.15 2.95 ;
        RECT  7.45 2.45 8.15 4.95 ;
        RECT  8.80 6.75 9.50 10.55 ;
        RECT  6.10 10.05 9.50 10.55 ;
        RECT  10.15 2.45 10.85 4.95 ;
        RECT  8.80 6.75 12.20 7.25 ;
        RECT  11.50 6.75 12.20 10.55 ;
        RECT  12.85 2.45 13.35 4.95 ;
        RECT  7.45 4.45 13.35 4.95 ;
        RECT  12.85 2.45 13.55 4.05 ;
    END
END EN2X3
MACRO EN2X4
    CLASS CORE ;
    FOREIGN EN2X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.70 6.75 5.40 10.55 ;
        RECT  4.80 3.45 5.50 5.10 ;
        RECT  4.80 4.60 8.20 5.10 ;
        RECT  7.50 3.40 8.20 7.25 ;
        RECT  7.25 4.60 8.20 7.25 ;
        RECT  8.90 6.75 9.60 9.60 ;
        RECT  4.70 6.75 12.30 7.25 ;
        RECT  11.60 6.75 12.30 9.60 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.10 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.10 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.35 7.20 4.05 11.00 ;
        RECT  6.05 7.70 6.75 11.00 ;
        RECT  14.45 7.70 15.15 11.00 ;
        RECT  17.15 7.70 17.85 11.00 ;
        RECT  19.85 7.15 20.55 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  10.20 2.00 10.90 4.00 ;
        RECT  12.90 2.00 13.60 4.00 ;
        RECT  15.60 2.00 16.30 4.00 ;
        RECT  18.30 2.00 19.00 4.00 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.90 3.60 1.40 6.05 ;
        RECT  0.90 3.60 1.65 4.30 ;
        RECT  1.85 5.55 2.35 10.55 ;
        RECT  1.85 7.45 2.55 8.15 ;
        RECT  1.85 9.85 2.55 10.55 ;
        RECT  0.90 5.55 4.60 6.05 ;
        RECT  3.45 2.45 4.15 4.15 ;
        RECT  3.90 5.55 4.60 6.25 ;
        RECT  6.15 2.45 6.85 4.15 ;
        RECT  7.55 7.70 8.25 10.55 ;
        RECT  3.45 2.45 9.55 2.95 ;
        RECT  8.85 2.45 9.55 4.95 ;
        RECT  10.25 7.70 10.95 10.55 ;
        RECT  11.55 2.45 12.25 4.95 ;
        RECT  12.95 6.75 13.65 10.55 ;
        RECT  7.55 10.05 13.65 10.55 ;
        RECT  14.25 2.45 14.95 4.95 ;
        RECT  15.80 6.75 16.50 10.55 ;
        RECT  16.95 2.45 17.65 4.95 ;
        RECT  12.95 6.75 19.20 7.25 ;
        RECT  18.50 6.75 19.20 10.55 ;
        RECT  19.65 2.45 20.15 4.95 ;
        RECT  8.85 4.45 20.15 4.95 ;
        RECT  19.65 2.45 20.35 4.05 ;
    END
END EN2X4
MACRO EN3X1
    CLASS CORE ;
    FOREIGN EN3X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.45 7.10 14.00 7.20 ;
        RECT  10.45 4.50 10.95 7.20 ;
        RECT  11.55 2.50 12.25 5.00 ;
        RECT  11.45 4.10 12.35 5.00 ;
        RECT  10.45 4.50 12.35 5.00 ;
        RECT  13.30 6.70 13.80 10.50 ;
        RECT  10.45 6.70 13.80 7.20 ;
        RECT  13.30 7.10 14.00 10.50 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.85 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.35 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.85 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  1.25 5.60 2.55 6.30 ;
        RECT  1.25 5.80 3.80 6.30 ;
        RECT  3.30 5.80 3.80 7.05 ;
        RECT  3.30 6.35 4.00 7.05 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.80 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.50 12.15 6.20 ;
        RECT  11.45 5.50 16.55 6.00 ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 7.50 3.50 11.00 ;
        RECT  5.50 8.85 6.20 11.00 ;
        RECT  11.80 7.75 12.80 8.45 ;
        RECT  12.30 7.75 12.80 11.00 ;
        RECT  15.65 7.10 16.35 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.35 2.00 3.05 3.90 ;
        RECT  6.90 2.00 7.60 3.85 ;
        RECT  14.30 2.00 15.00 3.90 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.25 4.40 0.75 10.45 ;
        RECT  0.25 7.55 1.15 10.45 ;
        RECT  0.75 2.70 1.50 4.90 ;
        RECT  3.55 2.50 4.00 5.10 ;
        RECT  3.30 4.40 4.00 5.10 ;
        RECT  3.55 2.50 4.05 4.90 ;
        RECT  0.25 4.40 4.05 4.90 ;
        RECT  4.15 7.85 4.85 10.45 ;
        RECT  4.55 3.50 5.05 7.35 ;
        RECT  4.55 3.50 5.25 4.20 ;
        RECT  3.55 2.50 6.25 3.00 ;
        RECT  5.75 2.50 6.25 4.90 ;
        RECT  4.15 7.85 7.70 8.35 ;
        RECT  5.75 4.35 7.75 4.90 ;
        RECT  7.00 7.85 7.70 10.45 ;
        RECT  7.25 4.35 7.75 6.35 ;
        RECT  7.25 5.65 7.95 6.35 ;
        RECT  4.55 6.85 8.95 7.35 ;
        RECT  8.25 4.35 8.95 5.05 ;
        RECT  8.45 4.35 8.95 10.45 ;
        RECT  8.35 6.85 8.95 10.45 ;
        RECT  8.35 8.45 9.05 10.45 ;
        RECT  9.80 3.20 9.95 8.20 ;
        RECT  9.45 3.40 9.95 8.20 ;
        RECT  9.45 7.70 10.75 8.20 ;
        RECT  9.80 3.20 10.50 3.90 ;
        RECT  9.45 3.40 10.50 3.90 ;
        RECT  10.05 7.70 10.75 10.50 ;
        RECT  10.05 9.30 11.80 10.00 ;
        RECT  12.90 2.50 13.60 4.10 ;
        RECT  13.10 2.50 13.60 4.90 ;
        RECT  15.65 2.50 16.15 4.90 ;
        RECT  13.10 4.40 16.15 4.90 ;
        RECT  15.65 2.50 16.35 4.10 ;
    END
END EN3X1
MACRO EN3X2
    CLASS CORE ;
    FOREIGN EN3X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  13.05 6.50 13.55 10.55 ;
        RECT  12.85 7.55 13.55 10.55 ;
        RECT  14.35 3.40 15.05 7.00 ;
        RECT  14.25 5.40 15.15 7.00 ;
        RECT  13.05 6.50 16.40 7.00 ;
        RECT  15.70 6.50 16.40 9.60 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.85 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.35 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.85 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  1.25 5.60 2.55 6.30 ;
        RECT  1.25 5.80 3.80 6.30 ;
        RECT  3.30 5.80 3.80 7.05 ;
        RECT  3.30 6.35 4.00 7.05 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 7.50 3.50 11.00 ;
        RECT  5.50 8.85 6.20 11.00 ;
        RECT  11.50 7.60 12.20 11.00 ;
        RECT  18.55 7.70 19.25 11.00 ;
        RECT  21.25 7.15 21.95 11.00 ;
        RECT  0.00 11.00 22.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.90 ;
        RECT  3.15 2.00 3.85 3.90 ;
        RECT  7.00 2.00 7.70 3.95 ;
        RECT  11.35 2.00 12.05 3.95 ;
        RECT  17.20 2.00 17.90 4.00 ;
        RECT  19.90 2.00 20.60 4.00 ;
        RECT  0.00 0.00 22.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.25 4.65 5.05 4.90 ;
        RECT  0.25 4.40 0.75 10.45 ;
        RECT  0.25 7.55 1.15 10.45 ;
        RECT  1.80 3.20 2.50 4.90 ;
        RECT  3.60 4.40 4.30 5.15 ;
        RECT  0.25 4.40 4.30 4.90 ;
        RECT  3.60 4.65 5.05 5.15 ;
        RECT  4.15 7.85 4.85 10.45 ;
        RECT  4.55 4.65 5.05 7.35 ;
        RECT  4.65 2.50 5.35 4.10 ;
        RECT  4.65 3.60 6.35 4.10 ;
        RECT  5.85 3.60 6.35 4.95 ;
        RECT  4.15 7.85 7.70 8.35 ;
        RECT  7.00 7.85 7.70 10.45 ;
        RECT  7.20 6.15 7.90 7.35 ;
        RECT  4.55 6.85 7.90 7.35 ;
        RECT  5.85 4.40 8.85 4.95 ;
        RECT  8.35 4.40 8.85 10.45 ;
        RECT  8.35 6.15 9.05 10.45 ;
        RECT  8.35 6.15 9.65 6.85 ;
        RECT  9.00 3.25 9.70 3.95 ;
        RECT  9.00 3.45 10.70 3.95 ;
        RECT  10.00 7.50 10.70 8.20 ;
        RECT  10.15 3.45 10.70 10.55 ;
        RECT  10.00 9.85 10.70 10.55 ;
        RECT  10.15 5.50 13.10 6.00 ;
        RECT  12.40 5.35 13.10 6.05 ;
        RECT  13.00 2.45 13.70 4.80 ;
        RECT  14.35 7.60 15.05 10.55 ;
        RECT  13.00 2.45 16.55 2.95 ;
        RECT  15.85 2.45 16.55 4.95 ;
        RECT  17.05 6.75 17.75 10.55 ;
        RECT  14.35 10.05 17.75 10.55 ;
        RECT  18.55 2.45 19.25 4.95 ;
        RECT  17.05 6.75 20.60 7.25 ;
        RECT  19.90 6.75 20.60 10.55 ;
        RECT  21.25 2.45 21.75 4.95 ;
        RECT  15.85 4.45 21.75 4.95 ;
        RECT  21.25 2.45 21.95 4.05 ;
    END
END EN3X2
MACRO EN3X3
    CLASS CORE ;
    FOREIGN EN3X3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  13.20 2.60 13.90 5.10 ;
        RECT  14.55 6.75 15.25 10.05 ;
        RECT  13.55 8.10 15.25 10.05 ;
        RECT  13.20 4.60 16.60 5.10 ;
        RECT  15.90 3.40 16.60 7.25 ;
        RECT  15.65 4.60 16.60 7.25 ;
        RECT  14.55 6.75 17.95 7.25 ;
        RECT  17.25 6.75 17.95 9.60 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.85 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.35 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.85 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  1.25 5.60 2.55 6.30 ;
        RECT  1.25 5.80 3.80 6.30 ;
        RECT  3.30 5.80 3.80 7.05 ;
        RECT  3.30 6.35 4.00 7.05 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 7.00 ;
        PORT
        LAYER M1M ;
        RECT  21.25 5.40 22.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 7.50 3.50 11.00 ;
        RECT  5.50 8.85 6.20 11.00 ;
        RECT  12.20 7.10 12.90 11.00 ;
        RECT  12.20 10.70 14.10 11.00 ;
        RECT  19.95 7.70 20.65 11.00 ;
        RECT  22.65 7.15 23.35 11.00 ;
        RECT  0.00 11.00 23.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.90 ;
        RECT  3.15 2.00 3.85 3.90 ;
        RECT  7.00 2.00 7.70 3.95 ;
        RECT  9.05 2.00 10.65 2.25 ;
        RECT  11.55 2.00 12.25 4.15 ;
        RECT  18.60 2.00 19.30 4.00 ;
        RECT  21.30 2.00 22.00 4.00 ;
        RECT  0.00 0.00 23.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.25 4.65 5.05 4.90 ;
        RECT  0.25 4.40 0.75 10.45 ;
        RECT  0.25 7.55 1.15 10.45 ;
        RECT  1.80 3.20 2.50 4.90 ;
        RECT  3.60 4.40 4.30 5.15 ;
        RECT  0.25 4.40 4.30 4.90 ;
        RECT  3.60 4.65 5.05 5.15 ;
        RECT  4.15 7.85 4.85 10.45 ;
        RECT  4.55 4.65 5.05 7.35 ;
        RECT  4.65 2.50 5.35 4.10 ;
        RECT  4.65 3.60 6.35 4.10 ;
        RECT  5.85 3.60 6.35 4.95 ;
        RECT  4.15 7.85 7.70 8.35 ;
        RECT  7.00 7.85 7.70 10.45 ;
        RECT  7.20 6.15 7.90 7.35 ;
        RECT  4.55 6.80 7.90 7.35 ;
        RECT  5.85 4.40 8.85 4.95 ;
        RECT  8.35 4.40 8.85 10.45 ;
        RECT  8.35 6.85 9.05 10.45 ;
        RECT  9.20 3.40 9.90 4.10 ;
        RECT  9.40 3.40 9.90 6.05 ;
        RECT  8.35 6.85 10.25 7.55 ;
        RECT  10.70 5.55 11.20 10.55 ;
        RECT  10.70 7.45 11.40 8.15 ;
        RECT  10.70 9.85 11.40 10.55 ;
        RECT  9.40 5.55 14.35 6.05 ;
        RECT  13.65 5.55 14.35 6.25 ;
        RECT  14.55 2.45 15.25 4.15 ;
        RECT  15.90 7.70 16.60 10.55 ;
        RECT  14.55 2.45 17.95 2.95 ;
        RECT  17.25 2.45 17.95 4.95 ;
        RECT  18.60 6.75 19.30 10.55 ;
        RECT  15.90 10.05 19.30 10.55 ;
        RECT  19.95 2.45 20.65 4.95 ;
        RECT  18.60 6.75 22.00 7.25 ;
        RECT  21.30 6.75 22.00 10.55 ;
        RECT  22.65 2.45 23.35 4.95 ;
        RECT  17.25 4.45 23.35 4.95 ;
    END
END EN3X3
MACRO EN3X4
    CLASS CORE ;
    FOREIGN EN3X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 29.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  13.10 6.75 13.80 10.55 ;
        RECT  13.20 3.45 13.90 5.10 ;
        RECT  13.20 4.60 16.60 5.10 ;
        RECT  15.90 3.40 16.60 7.25 ;
        RECT  15.65 4.60 16.60 7.25 ;
        RECT  17.30 6.75 18.00 9.60 ;
        RECT  13.10 6.75 20.70 7.25 ;
        RECT  20.00 6.75 20.70 9.60 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.85 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.85 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  1.25 5.60 2.55 6.30 ;
        RECT  1.25 5.80 3.80 6.30 ;
        RECT  3.30 5.80 3.80 7.05 ;
        RECT  3.30 6.35 4.00 7.05 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.10 ;
        PORT
        LAYER M1M ;
        RECT  24.05 5.40 24.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 7.50 3.50 11.00 ;
        RECT  5.50 8.85 6.20 11.00 ;
        RECT  11.75 7.20 12.45 11.00 ;
        RECT  14.45 7.70 15.15 11.00 ;
        RECT  22.85 7.70 23.55 11.00 ;
        RECT  25.55 7.70 26.25 11.00 ;
        RECT  28.25 7.15 28.95 11.00 ;
        RECT  0.00 11.00 29.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.90 ;
        RECT  3.15 2.00 3.85 3.90 ;
        RECT  7.00 2.00 7.70 3.95 ;
        RECT  8.95 2.00 10.55 2.50 ;
        RECT  18.60 2.00 19.30 4.10 ;
        RECT  21.30 2.00 22.00 4.10 ;
        RECT  24.00 2.00 24.70 4.00 ;
        RECT  26.70 2.00 27.40 4.00 ;
        RECT  0.00 0.00 29.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.25 4.65 5.05 4.90 ;
        RECT  0.25 4.40 0.75 10.45 ;
        RECT  0.25 7.55 1.15 10.45 ;
        RECT  1.80 3.20 2.50 4.90 ;
        RECT  3.60 4.40 4.30 5.15 ;
        RECT  0.25 4.40 4.30 4.90 ;
        RECT  3.60 4.65 5.05 5.15 ;
        RECT  4.15 7.85 4.85 10.45 ;
        RECT  4.55 4.65 5.05 7.30 ;
        RECT  4.65 2.50 5.35 4.10 ;
        RECT  4.65 3.60 6.35 4.10 ;
        RECT  5.85 3.60 6.35 4.95 ;
        RECT  4.15 7.85 7.70 8.35 ;
        RECT  7.00 7.85 7.70 10.45 ;
        RECT  7.20 6.15 7.90 7.30 ;
        RECT  4.55 6.80 7.90 7.30 ;
        RECT  5.85 4.40 8.85 4.95 ;
        RECT  8.35 4.40 8.85 10.45 ;
        RECT  8.35 7.35 9.05 10.45 ;
        RECT  8.35 4.95 9.80 5.65 ;
        RECT  9.50 3.50 10.20 4.20 ;
        RECT  9.50 3.70 11.05 4.20 ;
        RECT  10.25 7.45 11.05 8.15 ;
        RECT  10.55 3.70 11.05 10.55 ;
        RECT  10.25 9.85 11.05 10.55 ;
        RECT  11.85 2.45 12.55 4.15 ;
        RECT  12.30 5.55 13.00 6.25 ;
        RECT  10.55 5.75 13.00 6.25 ;
        RECT  14.55 2.45 15.25 4.15 ;
        RECT  15.95 7.70 16.65 10.55 ;
        RECT  11.85 2.45 17.95 2.95 ;
        RECT  17.25 2.45 17.95 5.05 ;
        RECT  18.65 7.70 19.35 10.55 ;
        RECT  19.95 2.55 20.65 5.05 ;
        RECT  21.35 6.75 22.05 10.55 ;
        RECT  15.95 10.05 22.05 10.55 ;
        RECT  22.65 2.55 23.35 5.05 ;
        RECT  17.25 4.55 23.35 5.05 ;
        RECT  24.20 6.75 24.90 10.55 ;
        RECT  25.35 2.45 26.05 4.95 ;
        RECT  21.35 6.75 27.60 7.25 ;
        RECT  26.90 6.75 27.60 10.55 ;
        RECT  22.65 4.45 28.55 4.95 ;
        RECT  28.05 2.45 28.55 4.95 ;
        RECT  17.25 4.55 28.55 4.95 ;
        RECT  28.05 2.45 28.75 4.05 ;
    END
END EN3X4
MACRO EO2X1
    CLASS CORE ;
    FOREIGN EO2X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  5.65 2.45 6.35 4.00 ;
        RECT  5.65 3.50 8.20 4.00 ;
        RECT  7.70 3.50 8.20 5.90 ;
        RECT  7.70 5.40 9.55 5.90 ;
        RECT  8.35 5.40 9.05 10.55 ;
        RECT  8.35 5.40 9.55 6.30 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.85 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.85 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 7.15 3.50 11.00 ;
        RECT  5.50 7.70 6.20 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 4.10 ;
        RECT  3.30 2.00 4.00 4.00 ;
        RECT  7.00 2.00 7.70 3.05 ;
        RECT  8.65 2.00 9.35 4.70 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 6.75 1.15 10.55 ;
        RECT  1.80 3.40 2.30 7.25 ;
        RECT  0.45 6.75 2.30 7.25 ;
        RECT  1.80 3.40 2.50 4.95 ;
        RECT  4.15 6.75 4.85 10.55 ;
        RECT  1.80 4.45 7.25 4.95 ;
        RECT  4.15 6.75 7.70 7.25 ;
        RECT  6.55 4.45 7.25 5.15 ;
        RECT  7.00 6.75 7.70 10.55 ;
    END
END EO2X1
MACRO EO2X2
    CLASS CORE ;
    FOREIGN EO2X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.65 3.40 9.35 5.00 ;
        RECT  11.45 2.45 12.20 5.00 ;
        RECT  11.70 2.45 12.20 9.60 ;
        RECT  11.50 7.10 12.20 9.60 ;
        RECT  11.45 4.10 12.35 5.00 ;
        RECT  8.65 4.50 12.35 5.00 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.95 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.95 ;
        PORT
        LAYER M1M ;
        RECT  2.55 5.60 3.25 6.30 ;
        RECT  7.25 5.40 8.15 6.30 ;
        RECT  2.55 5.80 8.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.10 7.70 3.80 11.00 ;
        RECT  5.80 8.65 6.50 11.00 ;
        RECT  8.50 8.65 9.20 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.10 2.00 3.80 4.05 ;
        RECT  5.80 2.00 6.50 4.00 ;
        RECT  12.85 2.00 13.55 4.05 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.60 6.75 1.30 10.55 ;
        RECT  1.40 2.55 2.10 4.15 ;
        RECT  1.60 2.55 2.10 7.25 ;
        RECT  4.45 2.45 5.15 4.95 ;
        RECT  4.45 7.70 5.15 10.55 ;
        RECT  7.15 7.70 7.85 10.55 ;
        RECT  7.30 2.45 8.00 4.95 ;
        RECT  4.45 4.45 8.00 4.95 ;
        RECT  9.05 6.20 9.55 7.25 ;
        RECT  0.60 6.75 9.55 7.25 ;
        RECT  7.30 2.45 10.70 2.95 ;
        RECT  4.45 7.70 10.85 8.20 ;
        RECT  10.00 2.45 10.70 4.05 ;
        RECT  10.15 7.15 10.85 10.55 ;
        RECT  10.55 6.00 11.25 6.70 ;
        RECT  9.05 6.20 11.25 6.70 ;
        RECT  12.85 7.15 13.55 10.55 ;
        RECT  10.15 10.05 13.55 10.55 ;
    END
END EO2X2
MACRO EO2X3
    CLASS CORE ;
    FOREIGN EO2X3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.70 3.40 9.40 5.00 ;
        RECT  11.40 2.50 12.10 5.00 ;
        RECT  14.50 3.15 14.95 9.60 ;
        RECT  14.25 3.15 14.95 5.00 ;
        RECT  14.50 4.10 15.00 9.60 ;
        RECT  14.30 7.10 15.00 9.60 ;
        RECT  14.25 4.10 15.15 5.00 ;
        RECT  8.70 4.50 15.15 5.00 ;
        RECT  14.50 6.20 17.70 6.70 ;
        RECT  17.00 6.20 17.70 10.55 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 8.05 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 8.05 ;
        PORT
        LAYER M1M ;
        RECT  2.75 5.60 3.45 6.30 ;
        RECT  7.25 5.40 8.15 6.30 ;
        RECT  2.75 5.80 8.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.10 7.70 3.80 11.00 ;
        RECT  5.80 8.65 6.50 11.00 ;
        RECT  8.50 8.65 9.20 11.00 ;
        RECT  11.20 8.65 11.90 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 4.15 ;
        RECT  3.30 2.00 4.00 4.05 ;
        RECT  6.00 2.00 6.70 4.00 ;
        RECT  12.90 2.00 13.60 3.85 ;
        RECT  15.60 2.00 16.30 3.85 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.60 6.75 1.30 10.55 ;
        RECT  1.80 3.45 2.30 7.25 ;
        RECT  1.80 3.45 2.50 4.15 ;
        RECT  4.45 7.70 5.15 10.55 ;
        RECT  4.65 2.45 5.35 4.95 ;
        RECT  7.15 7.70 7.85 10.55 ;
        RECT  7.35 2.45 8.05 4.95 ;
        RECT  4.65 4.45 8.05 4.95 ;
        RECT  7.35 2.45 10.75 2.95 ;
        RECT  9.85 7.70 10.55 10.55 ;
        RECT  10.05 2.45 10.75 4.05 ;
        RECT  11.65 6.20 12.15 7.25 ;
        RECT  0.60 6.75 12.15 7.25 ;
        RECT  4.45 7.70 13.65 8.20 ;
        RECT  12.95 7.15 13.65 10.55 ;
        RECT  13.35 6.00 14.05 6.70 ;
        RECT  11.65 6.20 14.05 6.70 ;
        RECT  15.65 7.15 16.35 10.55 ;
        RECT  12.95 10.05 16.35 10.55 ;
    END
END EO2X3
MACRO EO2X4
    CLASS CORE ;
    FOREIGN EO2X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.55 3.40 12.25 5.00 ;
        RECT  14.25 3.40 14.95 5.00 ;
        RECT  16.95 6.20 17.45 9.60 ;
        RECT  16.75 7.10 17.45 9.60 ;
        RECT  18.45 2.45 18.95 6.70 ;
        RECT  18.45 2.45 19.15 5.00 ;
        RECT  18.45 4.10 19.35 5.00 ;
        RECT  11.55 4.50 19.35 5.00 ;
        RECT  16.95 6.20 20.15 6.70 ;
        RECT  19.45 6.20 20.15 9.60 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 10.15 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 10.15 ;
        PORT
        LAYER M1M ;
        RECT  2.75 5.60 3.45 6.30 ;
        RECT  10.05 5.40 10.95 6.30 ;
        RECT  2.75 5.80 10.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.10 7.70 3.80 11.00 ;
        RECT  5.80 8.65 6.50 11.00 ;
        RECT  8.50 8.65 9.20 11.00 ;
        RECT  11.20 8.65 11.90 11.00 ;
        RECT  13.90 8.65 14.60 11.00 ;
        RECT  0.00 11.00 22.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 4.15 ;
        RECT  3.30 2.00 4.00 4.05 ;
        RECT  6.00 2.00 6.70 4.00 ;
        RECT  8.70 2.00 9.40 4.00 ;
        RECT  17.10 2.00 17.80 4.05 ;
        RECT  19.80 2.00 20.50 4.05 ;
        RECT  0.00 0.00 22.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.60 6.75 1.30 10.55 ;
        RECT  1.80 3.45 2.30 7.25 ;
        RECT  1.80 3.45 2.50 4.15 ;
        RECT  4.45 7.70 5.15 10.55 ;
        RECT  4.65 2.45 5.35 4.95 ;
        RECT  7.15 7.70 7.85 10.55 ;
        RECT  7.35 2.45 8.05 4.95 ;
        RECT  9.85 7.70 10.55 10.55 ;
        RECT  10.20 2.45 10.90 4.95 ;
        RECT  4.65 4.45 10.90 4.95 ;
        RECT  12.55 7.70 13.25 10.55 ;
        RECT  12.90 2.45 13.60 4.05 ;
        RECT  13.95 6.20 14.45 7.25 ;
        RECT  0.60 6.75 14.45 7.25 ;
        RECT  4.45 7.70 16.10 8.20 ;
        RECT  10.20 2.45 16.30 2.95 ;
        RECT  15.40 7.15 16.10 10.55 ;
        RECT  15.60 2.45 16.30 4.05 ;
        RECT  15.80 6.00 16.50 6.70 ;
        RECT  13.95 6.20 16.50 6.70 ;
        RECT  18.10 7.15 18.80 10.55 ;
        RECT  20.80 7.15 21.50 10.55 ;
        RECT  15.40 10.05 21.50 10.55 ;
    END
END EO2X4
MACRO EO3X1
    CLASS CORE ;
    FOREIGN EO3X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  14.90 3.55 15.60 4.25 ;
        RECT  15.10 3.55 15.60 6.00 ;
        RECT  15.10 5.50 19.35 6.00 ;
        RECT  18.35 5.40 18.45 10.50 ;
        RECT  17.75 5.50 18.45 10.50 ;
        RECT  18.35 5.40 19.35 6.30 ;
        RECT  17.75 5.50 19.35 6.30 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.85 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.85 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.35 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.85 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.45 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 7.10 3.50 11.00 ;
        RECT  5.50 8.15 6.20 11.00 ;
        RECT  12.20 7.10 12.90 11.00 ;
        RECT  14.90 7.50 15.60 11.00 ;
        RECT  0.00 11.00 19.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.85 ;
        RECT  3.15 2.00 3.85 3.85 ;
        RECT  7.85 2.00 8.55 4.45 ;
        RECT  9.85 2.00 10.55 3.85 ;
        RECT  12.55 2.00 13.25 3.85 ;
        RECT  17.10 2.00 17.80 3.80 ;
        RECT  0.00 0.00 19.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 4.35 0.95 10.50 ;
        RECT  0.45 7.10 1.15 10.50 ;
        RECT  1.80 3.15 2.50 4.85 ;
        RECT  4.35 2.55 4.85 4.85 ;
        RECT  0.45 4.35 4.85 4.85 ;
        RECT  4.15 7.10 4.85 10.50 ;
        RECT  5.50 3.80 6.35 4.50 ;
        RECT  5.85 3.80 6.35 6.65 ;
        RECT  4.35 2.55 7.35 3.05 ;
        RECT  4.15 7.10 7.70 7.65 ;
        RECT  6.85 2.55 7.35 5.65 ;
        RECT  6.85 4.95 7.55 5.65 ;
        RECT  7.00 7.10 7.70 10.50 ;
        RECT  8.15 4.95 8.85 6.65 ;
        RECT  5.85 6.15 8.85 6.65 ;
        RECT  8.35 4.95 8.85 10.50 ;
        RECT  8.35 7.10 9.05 10.50 ;
        RECT  10.05 4.35 10.55 10.50 ;
        RECT  9.85 7.10 10.55 10.50 ;
        RECT  11.20 3.15 11.90 4.85 ;
        RECT  13.75 2.55 14.25 4.85 ;
        RECT  10.05 4.35 14.25 4.85 ;
        RECT  13.75 6.50 14.25 10.50 ;
        RECT  13.55 7.10 14.25 10.50 ;
        RECT  13.75 2.55 16.60 3.05 ;
        RECT  13.75 6.50 16.90 7.00 ;
        RECT  16.10 2.55 16.60 4.80 ;
        RECT  16.10 4.30 17.55 4.80 ;
        RECT  16.40 6.50 16.90 10.50 ;
        RECT  16.40 7.10 17.10 10.50 ;
        RECT  16.85 4.30 17.55 5.00 ;
    END
END EO3X1
MACRO EO3X2
    CLASS CORE ;
    FOREIGN EO3X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  18.45 3.40 19.15 5.00 ;
        RECT  21.25 2.45 22.00 5.00 ;
        RECT  21.50 2.45 22.00 9.60 ;
        RECT  21.30 7.10 22.00 9.60 ;
        RECT  21.25 4.10 22.15 5.00 ;
        RECT  18.45 4.50 22.15 5.00 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.85 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.85 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.35 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.95 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 7.10 3.50 11.00 ;
        RECT  5.50 8.15 6.20 11.00 ;
        RECT  12.90 7.70 13.60 11.00 ;
        RECT  15.60 8.65 16.30 11.00 ;
        RECT  18.30 8.65 19.00 11.00 ;
        RECT  0.00 11.00 23.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.85 ;
        RECT  3.15 2.00 3.85 3.85 ;
        RECT  7.00 2.00 7.70 3.05 ;
        RECT  10.05 2.00 10.75 4.15 ;
        RECT  12.90 2.00 13.60 4.05 ;
        RECT  15.60 2.00 16.30 4.00 ;
        RECT  22.65 2.00 23.35 4.05 ;
        RECT  0.00 0.00 23.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 4.35 0.95 10.50 ;
        RECT  0.45 7.10 1.15 10.50 ;
        RECT  1.80 3.15 2.50 4.95 ;
        RECT  0.45 4.35 2.50 4.95 ;
        RECT  4.15 7.10 4.85 10.50 ;
        RECT  5.50 2.90 6.20 4.00 ;
        RECT  0.45 4.45 7.25 4.95 ;
        RECT  4.15 7.10 7.70 7.65 ;
        RECT  6.55 4.45 7.25 5.15 ;
        RECT  7.00 7.10 7.70 10.50 ;
        RECT  5.50 3.50 8.85 4.00 ;
        RECT  8.35 3.50 8.85 10.50 ;
        RECT  8.35 7.10 9.05 10.50 ;
        RECT  8.35 4.90 10.95 5.40 ;
        RECT  10.25 4.90 10.95 5.60 ;
        RECT  10.40 6.75 11.10 10.55 ;
        RECT  11.40 3.45 11.90 7.25 ;
        RECT  11.40 3.45 12.10 4.15 ;
        RECT  14.25 2.45 14.95 4.95 ;
        RECT  14.25 7.70 14.95 10.55 ;
        RECT  15.60 6.20 16.10 7.25 ;
        RECT  10.40 6.75 16.10 7.25 ;
        RECT  16.95 7.70 17.65 10.55 ;
        RECT  17.10 2.45 17.80 4.95 ;
        RECT  14.25 4.45 17.80 4.95 ;
        RECT  17.10 2.45 20.50 2.95 ;
        RECT  14.25 7.70 20.65 8.20 ;
        RECT  19.80 2.45 20.50 4.05 ;
        RECT  19.95 7.15 20.65 10.55 ;
        RECT  20.35 6.00 21.05 6.70 ;
        RECT  15.60 6.20 21.05 6.70 ;
        RECT  22.65 7.15 23.35 10.55 ;
        RECT  19.95 10.05 23.35 10.55 ;
    END
END EO3X2
MACRO EO3X3
    CLASS CORE ;
    FOREIGN EO3X3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 28.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  18.50 3.40 19.20 5.00 ;
        RECT  21.20 2.50 21.90 5.00 ;
        RECT  24.30 3.15 24.75 9.60 ;
        RECT  24.05 3.15 24.75 5.00 ;
        RECT  24.30 4.10 24.80 9.60 ;
        RECT  24.10 7.10 24.80 9.60 ;
        RECT  24.05 4.10 24.95 5.00 ;
        RECT  18.50 4.50 24.95 5.00 ;
        RECT  24.30 6.20 27.50 6.70 ;
        RECT  26.80 6.20 27.50 10.55 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.85 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.85 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.35 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 8.05 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 7.10 3.50 11.00 ;
        RECT  5.50 8.15 6.20 11.00 ;
        RECT  12.90 7.70 13.60 11.00 ;
        RECT  15.60 8.65 16.30 11.00 ;
        RECT  18.30 8.65 19.00 11.00 ;
        RECT  21.00 8.65 21.70 11.00 ;
        RECT  0.00 11.00 28.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.85 ;
        RECT  3.15 2.00 3.85 3.85 ;
        RECT  7.00 2.00 7.70 3.05 ;
        RECT  8.70 2.00 9.40 2.90 ;
        RECT  10.25 2.00 10.95 4.15 ;
        RECT  13.10 2.00 13.80 4.05 ;
        RECT  15.80 2.00 16.50 4.00 ;
        RECT  22.70 2.00 23.40 3.85 ;
        RECT  25.40 2.00 26.10 3.85 ;
        RECT  0.00 0.00 28.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 4.35 0.95 10.50 ;
        RECT  0.45 7.10 1.15 10.50 ;
        RECT  1.80 3.15 2.50 4.95 ;
        RECT  0.45 4.35 2.50 4.95 ;
        RECT  4.15 7.10 4.85 10.50 ;
        RECT  5.50 2.90 6.20 4.00 ;
        RECT  0.45 4.45 7.25 4.95 ;
        RECT  4.15 7.10 7.70 7.65 ;
        RECT  6.55 4.45 7.25 5.15 ;
        RECT  7.00 7.10 7.70 10.50 ;
        RECT  5.50 3.50 8.85 4.00 ;
        RECT  8.35 3.50 8.85 10.50 ;
        RECT  8.35 7.10 9.05 10.50 ;
        RECT  8.35 4.90 11.15 5.40 ;
        RECT  10.40 6.75 11.10 10.55 ;
        RECT  10.45 4.90 11.15 5.60 ;
        RECT  11.60 3.45 12.10 7.25 ;
        RECT  11.60 3.45 12.30 4.15 ;
        RECT  14.45 6.20 14.95 7.25 ;
        RECT  10.40 6.75 14.95 7.25 ;
        RECT  14.25 7.70 14.95 10.55 ;
        RECT  14.45 2.45 15.15 4.95 ;
        RECT  16.95 7.70 17.65 10.55 ;
        RECT  17.15 2.45 17.85 4.95 ;
        RECT  14.45 4.45 17.85 4.95 ;
        RECT  17.15 2.45 20.55 2.95 ;
        RECT  19.65 7.70 20.35 10.55 ;
        RECT  19.85 2.45 20.55 4.05 ;
        RECT  14.25 7.70 23.45 8.20 ;
        RECT  22.75 7.15 23.45 10.55 ;
        RECT  23.15 6.00 23.85 6.70 ;
        RECT  14.45 6.20 23.85 6.70 ;
        RECT  25.45 7.15 26.15 10.55 ;
        RECT  22.75 10.05 26.15 10.55 ;
    END
END EO3X3
MACRO EO3X4
    CLASS CORE ;
    FOREIGN EO3X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 32.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  21.35 3.40 22.05 5.00 ;
        RECT  24.05 3.40 24.75 5.00 ;
        RECT  26.75 6.20 27.25 9.60 ;
        RECT  26.55 7.10 27.25 9.60 ;
        RECT  28.25 2.45 28.75 6.70 ;
        RECT  28.25 2.45 28.95 5.00 ;
        RECT  28.25 4.10 29.15 5.00 ;
        RECT  21.35 4.50 29.15 5.00 ;
        RECT  26.75 6.20 29.95 6.70 ;
        RECT  29.25 6.20 29.95 9.60 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.85 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.85 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.35 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 10.15 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 7.10 3.50 11.00 ;
        RECT  5.50 8.15 6.20 11.00 ;
        RECT  12.90 7.70 13.60 11.00 ;
        RECT  15.60 8.65 16.30 11.00 ;
        RECT  18.30 8.65 19.00 11.00 ;
        RECT  21.00 8.65 21.70 11.00 ;
        RECT  23.70 8.65 24.40 11.00 ;
        RECT  0.00 11.00 32.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.85 ;
        RECT  3.15 2.00 3.85 3.85 ;
        RECT  7.00 2.00 7.70 3.05 ;
        RECT  8.70 2.00 9.40 2.90 ;
        RECT  10.25 2.00 10.95 4.15 ;
        RECT  13.10 2.00 13.80 4.05 ;
        RECT  15.80 2.00 16.50 4.00 ;
        RECT  18.50 2.00 19.20 4.00 ;
        RECT  26.90 2.00 27.60 4.05 ;
        RECT  29.60 2.00 30.30 4.05 ;
        RECT  0.00 0.00 32.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 4.35 0.95 10.50 ;
        RECT  0.45 7.10 1.15 10.50 ;
        RECT  1.80 3.15 2.50 4.95 ;
        RECT  0.45 4.35 2.50 4.95 ;
        RECT  4.15 7.10 4.85 10.50 ;
        RECT  5.50 2.90 6.20 4.00 ;
        RECT  0.45 4.45 7.25 4.95 ;
        RECT  4.15 7.10 7.70 7.65 ;
        RECT  6.55 4.45 7.25 5.15 ;
        RECT  7.00 7.10 7.70 10.50 ;
        RECT  5.50 3.50 8.85 4.00 ;
        RECT  8.35 3.50 8.85 10.50 ;
        RECT  8.35 7.10 9.05 10.50 ;
        RECT  8.35 4.90 11.15 5.40 ;
        RECT  10.40 6.75 11.10 10.55 ;
        RECT  10.45 4.90 11.15 5.60 ;
        RECT  11.60 3.45 12.10 7.25 ;
        RECT  11.60 3.45 12.30 4.15 ;
        RECT  14.25 7.70 14.95 10.55 ;
        RECT  14.45 2.45 15.15 4.95 ;
        RECT  14.75 6.20 15.25 7.25 ;
        RECT  10.40 6.75 15.25 7.25 ;
        RECT  16.95 7.70 17.65 10.55 ;
        RECT  17.15 2.45 17.85 4.95 ;
        RECT  19.65 7.70 20.35 10.55 ;
        RECT  20.00 2.45 20.70 4.95 ;
        RECT  14.45 4.45 20.70 4.95 ;
        RECT  22.35 7.70 23.05 10.55 ;
        RECT  22.70 2.45 23.40 4.05 ;
        RECT  14.25 7.70 25.90 8.20 ;
        RECT  20.00 2.45 26.10 2.95 ;
        RECT  25.20 7.15 25.90 10.55 ;
        RECT  25.40 2.45 26.10 4.05 ;
        RECT  25.60 6.00 26.30 6.70 ;
        RECT  14.75 6.20 26.30 6.70 ;
        RECT  27.90 7.15 28.60 10.55 ;
        RECT  30.60 7.15 31.30 10.55 ;
        RECT  25.20 10.05 31.30 10.55 ;
    END
END EO3X4
MACRO FAX1
    CLASS CORE ;
    FOREIGN FAX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 25.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.65 6.30 ;
        RECT  1.15 3.75 1.65 9.60 ;
        RECT  1.15 3.75 1.90 4.45 ;
        RECT  1.15 7.90 1.90 9.60 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M2M ;
        RECT  18.50 4.00 19.10 8.85 ;
        RECT  18.50 4.00 19.30 5.10 ;
        RECT  18.50 8.05 19.30 8.85 ;
        LAYER M1M ;
        RECT  18.45 3.75 19.35 5.00 ;
        RECT  18.45 8.00 19.35 9.65 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  24.05 6.70 24.95 7.60 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.20 ;
        PORT
        LAYER M1M ;
        RECT  14.25 6.70 15.50 7.60 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.20 ;
        PORT
        LAYER M1M ;
        RECT  7.15 5.40 8.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.55 7.90 3.25 11.00 ;
        RECT  5.40 9.85 6.10 11.00 ;
        RECT  8.10 9.85 8.80 11.00 ;
        RECT  14.45 8.05 15.15 11.00 ;
        RECT  17.15 8.05 17.85 11.00 ;
        RECT  20.35 8.05 21.05 11.00 ;
        RECT  0.00 11.00 25.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.55 2.00 3.25 4.45 ;
        RECT  7.50 2.00 8.20 4.45 ;
        RECT  10.20 2.00 10.90 4.45 ;
        RECT  17.15 2.00 17.85 4.45 ;
        RECT  21.35 2.00 22.05 4.35 ;
        RECT  0.00 0.00 25.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.10 6.75 2.80 7.45 ;
        RECT  4.15 3.75 4.85 4.45 ;
        RECT  4.05 8.85 4.75 10.55 ;
        RECT  4.35 3.75 4.85 7.25 ;
        RECT  4.60 7.70 5.30 8.40 ;
        RECT  6.75 8.85 7.45 10.55 ;
        RECT  8.85 3.80 9.55 5.40 ;
        RECT  4.05 8.85 11.10 9.35 ;
        RECT  10.60 8.85 11.10 10.55 ;
        RECT  10.80 7.70 11.50 8.40 ;
        RECT  4.60 7.90 11.50 8.40 ;
        RECT  11.55 3.75 12.25 5.40 ;
        RECT  8.85 4.90 12.25 5.40 ;
        RECT  11.95 6.75 12.45 9.55 ;
        RECT  11.55 8.85 12.45 9.55 ;
        RECT  12.90 3.75 13.40 7.25 ;
        RECT  2.10 6.75 13.40 7.25 ;
        RECT  12.90 3.75 13.60 4.45 ;
        RECT  12.90 8.85 13.60 10.55 ;
        RECT  10.60 10.05 13.60 10.55 ;
        RECT  14.80 3.75 15.50 6.25 ;
        RECT  14.10 5.55 15.50 6.25 ;
        RECT  16.00 6.95 16.50 9.65 ;
        RECT  15.80 8.05 16.50 9.65 ;
        RECT  18.05 5.75 18.75 6.45 ;
        RECT  20.00 3.70 20.70 5.30 ;
        RECT  16.00 6.95 22.20 7.45 ;
        RECT  21.70 6.95 22.20 10.55 ;
        RECT  22.70 5.75 23.20 9.60 ;
        RECT  22.70 3.70 23.40 5.30 ;
        RECT  20.00 4.80 23.40 5.30 ;
        RECT  22.70 8.00 23.40 9.60 ;
        RECT  24.05 3.70 24.55 6.25 ;
        RECT  14.10 5.75 24.55 6.25 ;
        RECT  24.05 3.70 24.75 4.40 ;
        RECT  24.05 8.05 24.75 10.55 ;
        RECT  21.70 10.05 24.75 10.55 ;
        LAYER V1M ;
        RECT  18.40 7.95 19.40 8.95 ;
        RECT  18.40 4.05 19.40 5.05 ;
    END
END FAX1
MACRO FAX2
    CLASS CORE ;
    FOREIGN FAX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 25.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.65 6.30 ;
        RECT  1.15 2.70 1.65 10.50 ;
        RECT  1.15 2.70 1.90 4.50 ;
        RECT  1.15 7.10 1.90 10.50 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M2M ;
        RECT  18.50 4.00 19.30 5.10 ;
        RECT  18.70 4.00 19.30 8.60 ;
        RECT  18.60 7.80 19.40 8.60 ;
        LAYER M1M ;
        RECT  18.55 7.75 19.45 8.65 ;
        RECT  18.45 2.70 19.20 5.00 ;
        RECT  18.45 4.10 19.35 5.00 ;
        RECT  18.70 7.75 19.45 10.50 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  24.05 6.70 24.95 7.60 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.20 ;
        PORT
        LAYER M1M ;
        RECT  14.25 6.70 15.50 7.60 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.20 ;
        PORT
        LAYER M1M ;
        RECT  7.15 5.40 8.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.55 7.10 3.25 11.00 ;
        RECT  5.40 9.85 6.10 11.00 ;
        RECT  8.10 9.85 8.80 11.00 ;
        RECT  14.45 8.05 15.15 11.00 ;
        RECT  17.35 7.75 18.05 11.00 ;
        RECT  20.35 8.05 21.05 11.00 ;
        RECT  0.00 11.00 25.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.55 2.00 3.25 4.50 ;
        RECT  7.50 2.00 8.20 4.45 ;
        RECT  10.20 2.00 10.90 4.45 ;
        RECT  17.15 2.00 17.85 4.50 ;
        RECT  21.35 2.00 22.05 4.35 ;
        RECT  0.00 0.00 25.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.10 5.45 2.80 6.15 ;
        RECT  4.15 3.75 4.85 4.45 ;
        RECT  2.10 5.45 4.85 5.95 ;
        RECT  4.05 8.85 4.75 10.55 ;
        RECT  4.35 3.75 4.85 7.25 ;
        RECT  4.60 7.70 5.30 8.40 ;
        RECT  6.75 8.85 7.45 10.55 ;
        RECT  8.85 3.80 9.55 5.40 ;
        RECT  4.05 8.85 11.10 9.35 ;
        RECT  10.60 8.85 11.10 10.55 ;
        RECT  10.80 7.70 11.50 8.40 ;
        RECT  4.60 7.90 11.50 8.40 ;
        RECT  11.55 3.75 12.25 5.40 ;
        RECT  8.85 4.90 12.25 5.40 ;
        RECT  11.95 6.75 12.45 9.55 ;
        RECT  11.55 8.85 12.45 9.55 ;
        RECT  12.90 3.75 13.40 7.25 ;
        RECT  4.35 6.75 13.40 7.25 ;
        RECT  12.90 3.75 13.60 4.45 ;
        RECT  12.90 8.85 13.60 10.55 ;
        RECT  10.60 10.05 13.60 10.55 ;
        RECT  14.65 3.75 15.35 6.25 ;
        RECT  14.30 5.55 15.35 6.25 ;
        RECT  16.00 6.75 16.50 9.65 ;
        RECT  15.80 8.05 16.50 9.65 ;
        RECT  18.05 5.55 18.75 6.25 ;
        RECT  20.00 3.70 20.70 5.30 ;
        RECT  16.00 6.75 22.20 7.25 ;
        RECT  21.70 6.75 22.20 10.55 ;
        RECT  22.70 5.75 23.20 9.60 ;
        RECT  22.70 3.70 23.40 5.30 ;
        RECT  20.00 4.80 23.40 5.30 ;
        RECT  22.70 8.00 23.40 9.60 ;
        RECT  24.05 3.70 24.55 6.25 ;
        RECT  14.30 5.75 24.55 6.25 ;
        RECT  24.05 3.70 24.75 4.40 ;
        RECT  24.05 8.05 24.75 10.55 ;
        RECT  21.70 10.05 24.75 10.55 ;
        LAYER V1M ;
        RECT  18.40 4.05 19.40 5.05 ;
        RECT  18.40 7.95 19.40 8.95 ;
    END
END FAX2

MACRO FAX3
    CLASS CORE ;
    FOREIGN FAX3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 26.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.80 3.40 2.55 4.15 ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  2.05 3.40 2.55 9.80 ;
        RECT  1.80 7.10 2.55 9.80 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M2M ;
        RECT  18.50 4.00 19.30 5.10 ;
        RECT  18.70 4.00 19.30 8.60 ;
        RECT  18.50 7.80 19.30 8.60 ;
        LAYER M1M ;
        RECT  18.45 7.75 19.80 8.65 ;
        RECT  18.60 3.70 19.35 5.00 ;
        RECT  18.45 4.10 19.35 5.00 ;
        RECT  19.10 7.75 19.80 10.50 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  25.45 6.70 26.35 7.60 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.20 ;
        PORT
        LAYER M1M ;
        RECT  14.25 6.70 15.15 7.60 ;
        RECT  14.25 6.85 15.95 7.60 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.20 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.25 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.10 1.15 11.00 ;
        RECT  3.15 7.10 3.85 11.00 ;
        RECT  6.00 9.85 6.70 11.00 ;
        RECT  8.70 9.85 9.40 11.00 ;
        RECT  14.90 8.05 15.60 11.00 ;
        RECT  17.75 9.15 18.45 11.00 ;
        RECT  20.45 8.05 22.45 11.00 ;
        RECT  0.00 11.00 26.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 4.15 ;
        RECT  3.15 2.00 3.85 4.15 ;
        RECT  8.00 2.00 8.70 4.45 ;
        RECT  10.70 2.00 11.40 4.45 ;
        RECT  17.25 2.00 17.95 4.40 ;
        RECT  19.95 2.00 20.65 4.40 ;
        RECT  23.00 2.00 23.70 2.85 ;
        RECT  0.00 0.00 26.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.05 5.45 3.75 6.15 ;
        RECT  4.65 3.75 5.35 4.45 ;
        RECT  3.05 5.45 5.35 5.95 ;
        RECT  4.85 3.75 5.35 7.25 ;
        RECT  4.65 8.85 5.35 10.50 ;
        RECT  5.10 7.70 5.80 8.40 ;
        RECT  7.35 8.85 8.05 10.50 ;
        RECT  8.75 5.85 9.30 7.25 ;
        RECT  4.85 6.75 9.30 7.25 ;
        RECT  9.35 3.80 10.05 5.40 ;
        RECT  4.65 8.85 11.55 9.35 ;
        RECT  11.05 8.85 11.55 10.50 ;
        RECT  11.40 6.80 11.90 8.20 ;
        RECT  5.10 7.70 11.90 8.20 ;
        RECT  11.40 6.80 12.10 7.50 ;
        RECT  12.40 7.95 12.90 9.50 ;
        RECT  12.05 3.75 12.75 5.40 ;
        RECT  9.35 4.90 12.75 5.40 ;
        RECT  12.65 5.85 12.90 9.50 ;
        RECT  12.05 8.80 12.90 9.50 ;
        RECT  12.65 5.85 13.15 8.45 ;
        RECT  12.40 7.95 13.15 8.45 ;
        RECT  13.40 3.75 13.90 6.35 ;
        RECT  8.75 5.85 13.90 6.35 ;
        RECT  13.40 3.75 14.10 4.45 ;
        RECT  13.40 8.85 14.10 10.50 ;
        RECT  11.05 10.00 14.10 10.50 ;
        RECT  14.90 3.75 15.60 6.25 ;
        RECT  14.40 5.55 15.60 6.25 ;
        RECT  16.45 6.75 16.95 9.65 ;
        RECT  16.25 8.05 16.95 9.65 ;
        RECT  18.15 5.55 18.85 6.25 ;
        RECT  21.50 3.70 22.20 4.45 ;
        RECT  16.45 6.75 23.60 7.25 ;
        RECT  23.10 6.75 23.60 10.55 ;
        RECT  24.10 5.75 24.60 9.60 ;
        RECT  24.10 3.70 24.80 4.45 ;
        RECT  21.50 3.95 24.80 4.45 ;
        RECT  24.10 8.00 24.80 9.60 ;
        RECT  25.45 3.70 25.95 6.25 ;
        RECT  14.40 5.75 25.95 6.25 ;
        RECT  25.45 3.70 26.15 4.40 ;
        RECT  25.45 8.05 26.15 10.55 ;
        RECT  23.10 10.05 26.15 10.55 ;
        LAYER V1M ;
        RECT  18.40 7.95 19.40 8.95 ;
        RECT  18.40 4.05 19.40 5.05 ;
    END
END FAX3
MACRO FAX3_YA_SIRENEVIY_TUMAN
    CLASS CORE ;
    FOREIGN FAX3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 26.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.80 3.40 2.55 4.15 ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  2.05 3.40 2.55 9.80 ;
        RECT  1.80 7.10 2.55 9.80 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M2M ;
        RECT  18.50 4.00 19.30 5.10 ;
        RECT  18.70 4.00 19.30 8.60 ;
        RECT  18.50 7.80 19.30 8.60 ;
        LAYER M1M ;
        RECT  18.45 7.75 19.80 8.65 ;
        RECT  18.60 3.70 19.35 5.00 ;
        RECT  18.45 4.10 19.35 5.00 ;
        RECT  19.10 7.75 19.80 10.50 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  25.45 6.70 26.35 7.60 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.20 ;
        PORT
        LAYER M1M ;
        RECT  14.25 6.70 15.15 7.60 ;
        RECT  14.25 6.85 15.95 7.60 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.20 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.25 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.10 1.15 11.00 ;
        RECT  3.15 7.10 3.85 11.00 ;
        RECT  6.00 9.85 6.70 11.00 ;
        RECT  8.70 9.85 9.40 11.00 ;
        RECT  14.90 8.05 15.60 11.00 ;
        RECT  17.75 9.15 18.45 11.00 ;
        RECT  20.45 8.05 22.45 11.00 ;
        RECT  0.00 11.00 26.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 4.15 ;
        RECT  3.15 2.00 3.85 4.15 ;
        RECT  8.00 2.00 8.70 4.45 ;
        RECT  10.70 2.00 11.40 4.45 ;
        RECT  17.25 2.00 17.95 4.40 ;
        RECT  19.95 2.00 20.65 4.40 ;
        RECT  23.00 2.00 23.70 2.85 ;
        RECT  0.00 0.00 26.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.05 5.45 3.75 6.15 ;
        RECT  4.65 3.75 5.35 4.45 ;
        RECT  3.05 5.45 5.35 5.95 ;
        RECT  4.85 3.75 5.35 7.25 ;
        RECT  4.65 8.85 5.35 10.50 ;
        RECT  5.10 7.70 5.80 8.40 ;
        RECT  7.35 8.85 8.05 10.50 ;
        RECT  8.75 5.85 9.30 7.25 ;
        RECT  4.85 6.75 9.30 7.25 ;
        RECT  9.35 3.80 10.05 5.40 ;
        RECT  4.65 8.85 11.55 9.35 ;
        RECT  11.05 8.85 11.55 10.50 ;
        RECT  11.40 6.80 11.90 8.20 ;
        RECT  5.10 7.70 11.90 8.20 ;
        RECT  11.40 6.80 12.10 7.50 ;
        RECT  12.40 7.95 12.90 9.50 ;
        RECT  12.05 3.75 12.75 5.40 ;
        RECT  9.35 4.90 12.75 5.40 ;
        RECT  12.65 5.85 12.90 9.50 ;
        RECT  12.05 8.80 12.90 9.50 ;
        RECT  12.65 5.85 13.15 8.45 ;
        RECT  12.40 7.95 13.15 8.45 ;
        RECT  13.40 3.75 13.90 6.35 ;
        RECT  8.75 5.85 13.90 6.35 ;
        RECT  13.40 3.75 14.10 4.45 ;
        RECT  13.40 8.85 14.10 10.50 ;
        RECT  11.05 10.00 14.10 10.50 ;
        RECT  14.90 3.75 15.60 6.25 ;
        RECT  14.40 5.55 15.60 6.25 ;
        RECT  16.45 6.75 16.95 9.65 ;
        RECT  16.25 8.05 16.95 9.65 ;
        RECT  18.15 5.55 18.85 6.25 ;
        RECT  21.50 3.70 22.20 4.45 ;
        RECT  16.45 6.75 23.60 7.25 ;
        RECT  23.10 6.75 23.60 10.55 ;
        RECT  24.10 5.75 24.60 9.60 ;
        RECT  24.10 3.70 24.80 4.45 ;
        RECT  21.50 3.95 24.80 4.45 ;
        RECT  24.10 8.00 24.80 9.60 ;
        RECT  25.45 3.70 25.95 6.25 ;
        RECT  14.40 5.75 25.95 6.25 ;
        RECT  25.45 3.70 26.15 4.40 ;
        RECT  25.45 8.05 26.15 10.55 ;
        RECT  23.10 10.05 26.15 10.55 ;
        LAYER V1M ;
        RECT  18.40 7.95 19.40 8.95 ;
        RECT  18.40 4.05 19.40 5.05 ;
    END
END FAX3
MACRO FAX4
    CLASS CORE ;
    FOREIGN FAX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 26.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.70 2.55 4.50 ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  2.05 2.70 2.55 10.50 ;
        RECT  1.80 7.10 2.55 10.50 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M2M ;
        RECT  18.50 4.00 19.30 5.10 ;
        RECT  18.70 4.00 19.30 8.60 ;
        RECT  18.50 7.80 19.30 8.60 ;
        LAYER M1M ;
        RECT  18.45 7.75 19.80 8.65 ;
        RECT  18.60 2.70 19.35 5.00 ;
        RECT  18.45 4.10 19.35 5.00 ;
        RECT  19.10 7.75 19.80 10.50 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  25.45 6.70 26.35 7.60 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.20 ;
        PORT
        LAYER M1M ;
        RECT  14.25 6.70 15.15 7.60 ;
        RECT  14.25 6.85 15.95 7.60 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.20 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.25 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.10 1.15 11.00 ;
        RECT  3.15 7.10 3.85 11.00 ;
        RECT  6.00 9.85 6.70 11.00 ;
        RECT  8.70 9.85 9.40 11.00 ;
        RECT  14.90 8.05 15.60 11.00 ;
        RECT  17.75 9.15 18.45 11.00 ;
        RECT  20.45 7.75 21.15 11.00 ;
        RECT  20.45 8.05 22.45 11.00 ;
        RECT  0.00 11.00 26.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 4.50 ;
        RECT  3.15 2.00 3.85 4.50 ;
        RECT  8.00 2.00 8.70 4.45 ;
        RECT  10.70 2.00 11.40 4.45 ;
        RECT  17.25 2.00 17.95 4.50 ;
        RECT  19.95 2.00 20.65 4.50 ;
        RECT  23.00 2.00 23.70 2.85 ;
        RECT  0.00 0.00 26.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.05 5.45 3.75 6.15 ;
        RECT  4.65 3.75 5.35 4.45 ;
        RECT  3.05 5.45 5.35 5.95 ;
        RECT  4.85 3.75 5.35 7.25 ;
        RECT  4.65 8.85 5.35 10.50 ;
        RECT  5.10 7.70 5.80 8.40 ;
        RECT  7.35 8.85 8.05 10.50 ;
        RECT  8.75 5.85 9.30 7.25 ;
        RECT  4.85 6.75 9.30 7.25 ;
        RECT  9.35 3.80 10.05 5.40 ;
        RECT  4.65 8.85 11.55 9.35 ;
        RECT  11.05 8.85 11.55 10.50 ;
        RECT  11.40 6.80 11.90 8.20 ;
        RECT  5.10 7.70 11.90 8.20 ;
        RECT  11.40 6.80 12.10 7.50 ;
        RECT  12.40 7.95 12.90 9.50 ;
        RECT  12.05 3.75 12.75 5.40 ;
        RECT  9.35 4.90 12.75 5.40 ;
        RECT  12.65 5.85 12.90 9.50 ;
        RECT  12.05 8.80 12.90 9.50 ;
        RECT  12.65 5.85 13.15 8.45 ;
        RECT  12.40 7.95 13.15 8.45 ;
        RECT  13.40 3.75 13.90 6.35 ;
        RECT  8.75 5.85 13.90 6.35 ;
        RECT  13.40 3.75 14.10 4.45 ;
        RECT  13.40 8.85 14.10 10.50 ;
        RECT  11.05 10.00 14.10 10.50 ;
        RECT  14.90 3.75 15.60 6.25 ;
        RECT  14.40 5.55 15.60 6.25 ;
        RECT  16.45 6.75 16.95 9.65 ;
        RECT  16.25 8.05 16.95 9.65 ;
        RECT  18.15 5.55 18.85 6.25 ;
        RECT  21.50 3.70 22.20 4.45 ;
        RECT  16.45 6.75 23.60 7.25 ;
        RECT  23.10 6.75 23.60 10.55 ;
        RECT  24.10 5.75 24.60 9.60 ;
        RECT  24.10 3.70 24.80 4.45 ;
        RECT  21.50 3.95 24.80 4.45 ;
        RECT  24.10 8.00 24.80 9.60 ;
        RECT  25.45 3.70 25.95 6.25 ;
        RECT  14.40 5.75 25.95 6.25 ;
        RECT  25.45 3.70 26.15 4.40 ;
        RECT  25.45 8.05 26.15 10.55 ;
        RECT  23.10 10.05 26.15 10.55 ;
        LAYER V1M ;
        RECT  18.40 7.95 19.40 8.95 ;
        RECT  18.40 4.05 19.40 5.05 ;
    END
END FAX4
MACRO FEED1
    CLASS CORE FEEDTHRU ;
    FOREIGN FEED1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 1.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.00 11.00 1.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.00 0.00 1.40 2.00 ;
        END
    END gnd!
END FEED1
MACRO FEED10
    CLASS CORE FEEDTHRU ;
    FOREIGN FEED10 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
END FEED10
MACRO FEED2
    CLASS CORE FEEDTHRU ;
    FOREIGN FEED2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.00 11.00 2.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.00 0.00 2.80 2.00 ;
        END
    END gnd!
END FEED2
MACRO FEED25
    CLASS CORE FEEDTHRU ;
    FOREIGN FEED25 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 35.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.00 11.00 35.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.00 0.00 35.00 2.00 ;
        END
    END gnd!
END FEED25
MACRO FEED5
    CLASS CORE FEEDTHRU ;
    FOREIGN FEED5 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.00 11.00 7.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.00 0.00 7.00 2.00 ;
        END
    END gnd!
END FEED5
MACRO HAX1
    CLASS CORE ;
    FOREIGN HAX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.25 2.45 10.75 9.15 ;
        RECT  10.05 7.45 10.75 9.15 ;
        RECT  9.90 2.45 10.95 3.70 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.25 2.45 1.20 3.70 ;
        RECT  0.70 2.45 1.20 9.10 ;
        RECT  0.50 7.45 1.20 9.10 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.05 9.30 3.95 10.20 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 7.50 2.55 11.00 ;
        RECT  4.70 7.50 5.40 11.00 ;
        RECT  0.45 10.65 5.40 11.00 ;
        RECT  8.55 7.70 9.25 11.00 ;
        RECT  10.05 10.10 10.75 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 2.00 2.55 3.15 ;
        RECT  7.05 4.05 7.75 4.75 ;
        RECT  8.55 2.00 9.05 4.55 ;
        RECT  7.05 4.05 9.05 4.55 ;
        RECT  8.55 2.00 9.25 3.15 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.65 6.35 2.35 7.05 ;
        RECT  3.35 2.45 3.85 8.15 ;
        RECT  3.35 6.55 4.05 8.15 ;
        RECT  4.35 4.05 5.05 4.75 ;
        RECT  3.35 2.45 4.90 3.15 ;
        RECT  4.55 4.05 5.05 5.80 ;
        RECT  5.05 6.35 5.75 7.05 ;
        RECT  1.65 6.55 5.75 7.05 ;
        RECT  4.55 5.30 6.70 5.80 ;
        RECT  5.90 2.65 6.40 4.75 ;
        RECT  5.70 4.05 6.40 4.75 ;
        RECT  6.20 5.30 6.70 10.55 ;
        RECT  6.20 6.75 6.90 10.55 ;
        RECT  7.20 2.45 7.90 3.15 ;
        RECT  5.90 2.65 7.90 3.15 ;
        RECT  9.10 6.35 9.60 7.25 ;
        RECT  6.20 6.75 9.60 7.25 ;
        RECT  9.10 6.35 9.80 7.05 ;
        RECT  6.20 6.75 9.80 7.05 ;
    END
END HAX1
MACRO HAX2
    CLASS CORE ;
    FOREIGN HAX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.05 2.45 10.75 4.20 ;
        RECT  10.25 2.45 10.75 10.55 ;
        RECT  10.05 7.45 10.75 10.55 ;
        RECT  10.05 2.45 10.95 3.70 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.25 2.45 1.15 3.70 ;
        RECT  0.45 2.45 0.95 10.50 ;
        RECT  0.45 2.45 1.15 4.15 ;
        RECT  0.45 7.10 1.15 10.50 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.05 9.30 3.95 10.20 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.10 2.50 11.00 ;
        RECT  4.70 7.50 5.40 11.00 ;
        RECT  8.60 7.70 9.30 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.15 ;
        RECT  7.05 4.05 7.75 4.75 ;
        RECT  8.70 2.00 9.40 4.55 ;
        RECT  7.05 4.05 9.40 4.55 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.45 6.55 5.75 6.60 ;
        RECT  1.45 5.90 2.15 6.60 ;
        RECT  3.35 2.45 3.85 8.15 ;
        RECT  1.45 6.10 3.85 6.60 ;
        RECT  3.35 6.55 4.05 8.15 ;
        RECT  4.35 4.10 5.05 4.80 ;
        RECT  3.35 2.45 5.00 3.15 ;
        RECT  4.55 4.10 5.05 5.80 ;
        RECT  5.05 6.35 5.75 7.05 ;
        RECT  3.35 6.55 5.75 7.05 ;
        RECT  4.55 5.30 6.70 5.80 ;
        RECT  5.90 2.65 6.40 4.75 ;
        RECT  5.70 4.05 6.40 4.75 ;
        RECT  6.20 5.30 6.70 10.55 ;
        RECT  6.20 6.75 6.90 10.55 ;
        RECT  7.20 2.45 7.90 3.15 ;
        RECT  5.90 2.65 7.90 3.15 ;
        RECT  9.10 6.35 9.60 7.25 ;
        RECT  6.20 6.75 9.60 7.25 ;
        RECT  9.10 6.35 9.80 7.05 ;
        RECT  6.20 6.75 9.80 7.05 ;
    END
END HAX2
MACRO HAX3
    CLASS CORE ;
    FOREIGN HAX3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.45 3.45 12.15 5.00 ;
        RECT  11.65 3.45 12.15 10.20 ;
        RECT  11.45 7.45 12.15 10.20 ;
        RECT  11.45 4.10 12.35 5.00 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.85 3.45 2.35 9.80 ;
        RECT  1.85 3.45 2.55 5.00 ;
        RECT  1.65 4.10 2.55 5.00 ;
        RECT  1.85 7.10 2.55 9.80 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  4.45 9.30 5.35 10.20 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.40 9.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 7.10 1.20 11.00 ;
        RECT  3.20 7.10 3.90 11.00 ;
        RECT  6.10 7.50 6.80 11.00 ;
        RECT  9.95 7.70 10.65 11.00 ;
        RECT  12.80 7.45 13.50 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 2.00 1.20 4.20 ;
        RECT  3.20 2.00 4.05 4.20 ;
        RECT  8.45 4.05 9.15 4.75 ;
        RECT  9.95 2.00 10.80 4.55 ;
        RECT  8.45 4.05 10.80 4.55 ;
        RECT  12.80 2.00 13.50 4.20 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.85 6.55 7.15 6.60 ;
        RECT  2.85 5.90 3.55 6.60 ;
        RECT  4.75 2.45 5.25 8.15 ;
        RECT  2.85 6.10 5.25 6.60 ;
        RECT  4.75 6.55 5.45 8.15 ;
        RECT  5.75 4.10 6.45 4.80 ;
        RECT  4.75 2.45 6.40 3.15 ;
        RECT  5.95 4.10 6.45 5.80 ;
        RECT  6.45 6.35 7.15 7.05 ;
        RECT  4.75 6.55 7.15 7.05 ;
        RECT  5.95 5.30 8.10 5.80 ;
        RECT  7.30 2.65 7.80 4.75 ;
        RECT  7.10 4.05 7.80 4.75 ;
        RECT  7.60 5.30 8.10 10.55 ;
        RECT  7.60 6.75 8.30 10.55 ;
        RECT  8.60 2.45 9.30 3.15 ;
        RECT  7.30 2.65 9.30 3.15 ;
        RECT  10.50 6.35 11.00 7.25 ;
        RECT  7.60 6.75 11.00 7.25 ;
        RECT  10.50 6.35 11.20 7.05 ;
        RECT  7.60 6.75 11.20 7.05 ;
    END
END HAX3
MACRO HAX4
    CLASS CORE ;
    FOREIGN HAX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.45 2.45 12.15 4.20 ;
        RECT  11.65 2.45 12.15 10.55 ;
        RECT  11.45 7.45 12.15 10.55 ;
        RECT  11.45 2.45 12.35 3.70 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.65 2.45 2.55 3.70 ;
        RECT  1.85 2.45 2.35 10.50 ;
        RECT  1.85 2.45 2.55 4.15 ;
        RECT  1.85 7.10 2.55 10.50 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  4.45 9.30 5.35 10.20 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.40 9.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 7.10 1.20 11.00 ;
        RECT  3.20 7.10 3.90 11.00 ;
        RECT  6.10 7.50 6.80 11.00 ;
        RECT  10.00 7.70 10.70 11.00 ;
        RECT  12.80 7.70 13.50 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 2.00 1.20 4.15 ;
        RECT  3.20 2.00 3.90 4.15 ;
        RECT  8.45 4.05 9.15 4.75 ;
        RECT  10.10 2.00 10.80 4.55 ;
        RECT  8.45 4.05 10.80 4.55 ;
        RECT  12.80 2.00 13.50 4.20 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.85 6.55 7.15 6.60 ;
        RECT  2.85 5.90 3.55 6.60 ;
        RECT  4.75 2.45 5.25 8.15 ;
        RECT  2.85 6.10 5.25 6.60 ;
        RECT  4.75 6.55 5.45 8.15 ;
        RECT  5.75 4.10 6.45 4.80 ;
        RECT  4.75 2.45 6.40 3.15 ;
        RECT  5.95 4.10 6.45 5.80 ;
        RECT  6.45 6.35 7.15 7.05 ;
        RECT  4.75 6.55 7.15 7.05 ;
        RECT  5.95 5.30 8.10 5.80 ;
        RECT  7.30 2.65 7.80 4.75 ;
        RECT  7.10 4.05 7.80 4.75 ;
        RECT  7.60 5.30 8.10 10.55 ;
        RECT  7.60 6.75 8.30 10.55 ;
        RECT  8.60 2.45 9.30 3.15 ;
        RECT  7.30 2.65 9.30 3.15 ;
        RECT  10.50 6.35 11.00 7.25 ;
        RECT  7.60 6.75 11.00 7.25 ;
        RECT  10.50 6.35 11.20 7.05 ;
        RECT  7.60 6.75 11.20 7.05 ;
    END
END HAX4
MACRO INCX12
    CLASS CORE ;
    FOREIGN INCX12 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.15 4.40 12.15 4.60 ;
        RECT  6.00 7.00 6.80 10.55 ;
        RECT  6.00 7.00 9.50 7.50 ;
        RECT  8.35 2.45 8.85 4.90 ;
        RECT  8.15 2.45 8.85 4.60 ;
        RECT  9.00 5.80 9.50 10.55 ;
        RECT  8.70 7.00 9.50 10.55 ;
        RECT  11.45 2.45 12.15 4.90 ;
        RECT  8.35 4.40 12.15 4.90 ;
        RECT  11.65 2.45 11.90 10.55 ;
        RECT  11.40 5.80 11.90 10.55 ;
        RECT  11.65 2.45 12.15 6.30 ;
        RECT  11.40 7.10 12.20 10.55 ;
        RECT  11.45 5.40 12.35 6.30 ;
        RECT  9.00 5.80 12.35 6.30 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.26 ;
        PORT
        LAYER M1M ;
        RECT  0.25 2.75 1.15 3.70 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 9.10 2.60 11.00 ;
        RECT  4.65 7.35 5.45 11.00 ;
        RECT  7.35 7.95 8.15 11.00 ;
        RECT  10.05 7.10 10.85 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.65 2.00 2.65 2.65 ;
        RECT  3.80 2.00 4.50 2.40 ;
        RECT  6.80 2.00 7.50 4.30 ;
        RECT  10.10 2.00 10.20 3.95 ;
        RECT  9.50 2.95 10.20 3.95 ;
        RECT  10.10 2.00 10.80 3.45 ;
        RECT  9.50 2.95 10.80 3.45 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.65 4.30 1.15 10.55 ;
        RECT  0.50 8.70 1.25 10.55 ;
        RECT  1.60 3.20 2.20 5.00 ;
        RECT  0.65 4.30 2.20 5.00 ;
        RECT  2.05 5.45 2.55 8.65 ;
        RECT  1.60 3.20 2.60 3.95 ;
        RECT  2.05 8.15 3.95 8.65 ;
        RECT  3.60 5.25 4.30 5.95 ;
        RECT  3.30 6.40 3.80 7.70 ;
        RECT  3.00 6.95 3.80 7.70 ;
        RECT  3.15 8.15 3.95 10.55 ;
        RECT  3.80 3.35 4.30 5.95 ;
        RECT  2.05 5.45 4.30 5.95 ;
        RECT  3.80 3.35 4.50 4.10 ;
        RECT  5.05 5.25 5.55 6.90 ;
        RECT  3.30 6.40 5.55 6.90 ;
        RECT  5.55 2.45 6.05 5.75 ;
        RECT  5.40 2.45 6.15 4.30 ;
        RECT  5.05 5.25 7.95 5.75 ;
        RECT  7.25 5.15 7.95 5.85 ;
    END
END INCX12
MACRO INCX16
    CLASS CORE ;
    FOREIGN INCX16 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.90 7.00 9.70 10.55 ;
        RECT  8.90 7.00 12.40 7.50 ;
        RECT  11.65 2.45 12.35 4.70 ;
        RECT  11.90 5.40 12.40 10.55 ;
        RECT  11.60 7.00 12.40 10.55 ;
        RECT  11.90 5.40 17.50 5.90 ;
        RECT  14.35 2.45 15.05 4.70 ;
        RECT  11.65 4.20 15.05 4.70 ;
        RECT  14.55 2.45 14.80 10.55 ;
        RECT  14.25 5.40 14.80 10.55 ;
        RECT  14.55 2.45 15.05 6.30 ;
        RECT  14.25 7.10 15.10 10.55 ;
        RECT  14.25 5.40 15.15 6.30 ;
        RECT  14.25 5.40 17.50 6.00 ;
        RECT  17.00 2.45 17.50 10.55 ;
        RECT  17.00 2.45 17.75 4.70 ;
        RECT  17.00 7.10 17.80 10.55 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.40 7.20 1.20 11.00 ;
        RECT  4.70 9.25 5.50 11.00 ;
        RECT  7.55 7.10 8.35 11.00 ;
        RECT  10.25 7.95 11.05 11.00 ;
        RECT  12.95 7.10 13.75 11.00 ;
        RECT  15.65 7.10 16.45 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.40 2.00 1.20 4.50 ;
        RECT  3.30 2.00 5.15 4.20 ;
        RECT  3.30 2.00 6.65 2.80 ;
        RECT  7.40 2.00 8.20 4.45 ;
        RECT  10.30 2.00 11.00 4.45 ;
        RECT  13.00 2.00 13.70 3.75 ;
        RECT  15.70 2.00 16.40 4.45 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.75 2.60 2.55 4.50 ;
        RECT  2.05 2.60 2.55 10.55 ;
        RECT  1.75 7.20 2.55 10.55 ;
        RECT  2.05 5.50 2.85 6.20 ;
        RECT  3.35 8.30 4.15 10.55 ;
        RECT  4.95 5.10 5.45 8.80 ;
        RECT  4.95 5.10 5.80 6.30 ;
        RECT  3.35 8.30 6.85 8.80 ;
        RECT  5.90 3.65 6.60 4.40 ;
        RECT  6.10 3.65 6.60 5.60 ;
        RECT  4.95 5.10 6.60 5.60 ;
        RECT  6.25 6.05 6.75 7.80 ;
        RECT  5.95 7.05 6.75 7.80 ;
        RECT  6.05 8.30 6.85 10.55 ;
        RECT  8.75 2.55 9.50 6.55 ;
        RECT  6.25 6.05 9.50 6.55 ;
        RECT  8.75 5.25 11.45 5.75 ;
        RECT  10.75 5.20 11.45 5.90 ;
    END
END INCX16
MACRO INCX20
    CLASS CORE ;
    FOREIGN INCX20 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.90 5.45 17.80 5.90 ;
        RECT  8.90 7.00 9.70 10.55 ;
        RECT  8.90 7.00 12.40 7.50 ;
        RECT  11.70 2.45 12.40 4.70 ;
        RECT  11.90 5.40 12.40 10.55 ;
        RECT  11.60 7.00 12.40 10.55 ;
        RECT  14.40 2.45 15.10 4.70 ;
        RECT  11.70 4.20 15.10 4.70 ;
        RECT  14.60 2.45 14.80 10.55 ;
        RECT  14.20 5.40 14.80 10.55 ;
        RECT  14.60 2.45 15.10 6.30 ;
        RECT  14.20 7.10 15.10 10.55 ;
        RECT  14.20 5.40 15.15 6.30 ;
        RECT  17.10 2.45 17.60 5.90 ;
        RECT  17.30 2.45 17.60 10.55 ;
        RECT  11.90 5.40 17.60 5.90 ;
        RECT  17.10 2.45 17.80 4.70 ;
        RECT  17.30 5.45 17.80 10.55 ;
        RECT  17.00 7.10 17.80 10.55 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.40 7.20 1.20 11.00 ;
        RECT  4.70 9.25 5.50 11.00 ;
        RECT  7.55 7.10 8.35 11.00 ;
        RECT  10.25 7.95 11.05 11.00 ;
        RECT  12.95 7.10 13.75 11.00 ;
        RECT  15.65 7.10 16.45 11.00 ;
        RECT  18.35 7.10 19.15 11.00 ;
        RECT  0.00 11.00 19.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.40 2.00 1.20 4.45 ;
        RECT  3.25 2.00 5.20 4.10 ;
        RECT  3.25 2.00 6.70 2.75 ;
        RECT  7.45 2.00 8.25 4.45 ;
        RECT  10.35 2.00 11.05 4.35 ;
        RECT  13.05 2.00 13.75 3.75 ;
        RECT  15.75 2.00 16.45 4.45 ;
        RECT  18.45 2.00 19.15 4.45 ;
        RECT  0.00 0.00 19.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.75 2.60 2.55 4.55 ;
        RECT  2.05 2.60 2.55 10.55 ;
        RECT  1.75 7.10 2.55 10.55 ;
        RECT  2.05 5.50 2.85 6.20 ;
        RECT  3.35 8.30 4.15 10.55 ;
        RECT  5.30 5.10 5.45 8.80 ;
        RECT  4.95 5.60 5.45 8.80 ;
        RECT  5.30 5.10 5.80 6.30 ;
        RECT  4.95 5.60 5.80 6.30 ;
        RECT  3.35 8.30 6.85 8.80 ;
        RECT  5.30 5.10 6.65 5.60 ;
        RECT  6.15 3.65 6.65 5.60 ;
        RECT  6.00 3.65 6.70 4.40 ;
        RECT  6.25 6.05 6.75 7.80 ;
        RECT  5.95 7.05 6.75 7.80 ;
        RECT  6.05 8.30 6.85 10.55 ;
        RECT  8.80 2.55 9.55 4.45 ;
        RECT  9.05 2.55 9.55 6.55 ;
        RECT  6.25 6.05 9.55 6.55 ;
        RECT  9.05 5.20 11.45 5.70 ;
        RECT  10.75 5.20 11.45 5.90 ;
    END
END INCX20
MACRO INCX3
    CLASS CORE ;
    FOREIGN INCX3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  5.85 7.10 7.95 7.95 ;
        RECT  7.25 2.45 7.95 4.60 ;
        RECT  7.45 2.45 7.95 10.55 ;
        RECT  7.15 7.10 7.95 10.55 ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.63 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.40 10.05 1.20 11.00 ;
        RECT  1.95 7.05 2.75 8.95 ;
        RECT  2.25 7.05 2.75 11.00 ;
        RECT  1.95 9.80 2.75 11.00 ;
        RECT  5.80 8.50 6.60 11.00 ;
        RECT  0.00 11.00 8.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.65 2.00 3.45 2.45 ;
        RECT  4.30 2.00 5.15 2.45 ;
        RECT  5.90 2.00 6.60 4.50 ;
        RECT  0.00 0.00 8.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.85 4.55 3.90 4.95 ;
        RECT  0.75 5.45 1.25 8.10 ;
        RECT  0.45 7.10 1.25 8.10 ;
        RECT  0.85 2.75 1.65 3.55 ;
        RECT  0.85 3.05 2.30 3.55 ;
        RECT  1.80 3.05 2.30 5.95 ;
        RECT  1.80 5.25 2.50 5.95 ;
        RECT  0.75 5.45 2.50 5.95 ;
        RECT  3.20 3.75 3.60 5.70 ;
        RECT  3.20 4.55 3.90 5.70 ;
        RECT  3.30 3.75 3.60 8.95 ;
        RECT  2.85 3.75 3.60 4.95 ;
        RECT  3.30 4.55 3.90 8.95 ;
        RECT  3.30 7.05 4.10 8.95 ;
        RECT  4.55 3.75 5.05 10.55 ;
        RECT  4.30 9.80 5.05 10.55 ;
        RECT  4.35 3.75 5.15 4.55 ;
        RECT  4.55 5.35 6.80 5.85 ;
        RECT  6.10 5.30 6.80 6.00 ;
    END
END INCX3
MACRO INCX4
    CLASS CORE ;
    FOREIGN INCX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  7.25 2.70 7.95 4.60 ;
        RECT  7.25 5.40 7.55 10.55 ;
        RECT  7.05 5.95 7.55 10.55 ;
        RECT  7.45 2.70 7.55 10.55 ;
        RECT  6.75 7.10 7.55 10.55 ;
        RECT  7.45 2.70 7.95 6.35 ;
        RECT  7.25 5.40 8.15 6.35 ;
        RECT  7.05 5.95 8.15 6.35 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.63 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.90 8.50 2.40 11.00 ;
        RECT  1.95 7.05 2.40 11.00 ;
        RECT  1.60 9.80 2.40 11.00 ;
        RECT  1.95 7.05 2.75 9.05 ;
        RECT  1.90 8.50 2.75 9.05 ;
        RECT  5.45 7.10 6.20 11.00 ;
        RECT  8.10 7.10 8.90 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.65 2.00 3.45 2.45 ;
        RECT  4.30 2.00 5.15 2.45 ;
        RECT  5.90 2.00 6.60 4.40 ;
        RECT  8.55 2.00 9.35 4.50 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.85 4.55 3.90 4.95 ;
        RECT  0.75 5.45 1.25 8.00 ;
        RECT  0.45 7.05 1.25 8.00 ;
        RECT  0.85 2.70 1.65 3.50 ;
        RECT  0.85 3.00 2.30 3.50 ;
        RECT  1.80 3.00 2.30 5.95 ;
        RECT  1.80 5.25 2.50 5.95 ;
        RECT  0.75 5.45 2.50 5.95 ;
        RECT  3.20 3.75 3.60 5.70 ;
        RECT  3.20 4.55 3.90 5.70 ;
        RECT  3.35 3.75 3.60 8.95 ;
        RECT  2.85 3.75 3.60 4.95 ;
        RECT  3.35 4.55 3.90 8.95 ;
        RECT  3.35 7.05 4.05 8.95 ;
        RECT  4.50 3.75 4.65 10.55 ;
        RECT  3.95 9.80 4.65 10.55 ;
        RECT  4.50 3.75 5.00 10.30 ;
        RECT  3.95 9.80 5.00 10.30 ;
        RECT  4.50 3.75 5.05 5.50 ;
        RECT  4.35 3.75 5.15 4.50 ;
        RECT  4.50 5.00 6.80 5.50 ;
        RECT  6.10 4.85 6.80 5.55 ;
    END
END INCX4
MACRO INCX8
    CLASS CORE ;
    FOREIGN INCX8 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  7.30 7.10 7.50 10.55 ;
        RECT  6.70 9.60 7.50 10.55 ;
        RECT  7.80 2.60 8.50 4.40 ;
        RECT  8.00 2.60 8.05 10.10 ;
        RECT  7.55 6.00 8.05 10.10 ;
        RECT  7.30 7.10 8.10 10.10 ;
        RECT  6.70 9.60 8.10 10.10 ;
        RECT  8.00 2.60 8.50 6.50 ;
        RECT  7.55 6.00 10.55 6.50 ;
        RECT  10.05 5.40 10.55 10.55 ;
        RECT  10.00 7.10 10.80 10.55 ;
        RECT  10.05 5.40 10.95 6.30 ;
        RECT  7.55 6.00 10.95 6.30 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.26 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.65 9.15 3.45 11.00 ;
        RECT  5.95 7.05 6.15 11.00 ;
        RECT  5.35 8.60 6.15 11.00 ;
        RECT  5.95 7.05 6.75 9.10 ;
        RECT  5.35 8.60 6.75 9.10 ;
        RECT  8.65 7.10 9.45 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.40 2.00 2.20 3.05 ;
        RECT  3.40 2.00 4.20 2.80 ;
        RECT  6.45 2.00 7.15 4.30 ;
        RECT  6.45 2.00 8.30 2.10 ;
        RECT  10.05 2.00 10.75 4.40 ;
        RECT  9.05 3.60 10.75 4.40 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.60 3.65 2.10 10.55 ;
        RECT  1.30 8.65 2.10 10.55 ;
        RECT  1.45 3.65 2.15 4.35 ;
        RECT  1.60 6.50 2.80 7.20 ;
        RECT  3.55 3.65 3.85 8.70 ;
        RECT  3.35 5.70 3.85 8.70 ;
        RECT  3.35 8.20 4.80 8.70 ;
        RECT  3.55 3.65 4.05 6.40 ;
        RECT  3.35 5.70 4.05 6.40 ;
        RECT  3.40 3.65 4.20 4.45 ;
        RECT  4.00 8.20 4.80 10.55 ;
        RECT  4.70 4.90 5.20 7.75 ;
        RECT  4.30 6.95 5.20 7.75 ;
        RECT  5.20 2.50 5.70 5.40 ;
        RECT  5.05 2.50 5.80 4.40 ;
        RECT  4.70 4.90 7.50 5.40 ;
        RECT  6.80 4.75 7.50 5.45 ;
    END
END INCX8
MACRO INX1
    CLASS CORE ;
    FOREIGN INX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M2M ;
        RECT  0.30 4.00 0.90 9.25 ;
        RECT  0.30 4.00 1.10 5.10 ;
        RECT  0.30 8.45 1.10 9.25 ;
        LAYER M1M ;
        RECT  0.25 3.80 1.15 5.00 ;
        RECT  0.25 8.40 1.60 9.30 ;
        RECT  0.25 3.80 1.75 4.50 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.90 7.10 2.55 7.80 ;
        RECT  2.05 7.10 2.55 11.00 ;
        RECT  0.90 9.80 2.55 11.00 ;
        RECT  0.00 11.00 2.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.05 2.00 1.75 3.15 ;
        RECT  0.00 0.00 2.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER V1M ;
        RECT  0.20 9.25 1.20 10.25 ;
        RECT  0.20 7.95 1.20 8.95 ;
        RECT  0.20 4.05 1.20 5.05 ;
    END
END INX1
MACRO INX12
    CLASS CORE ;
    FOREIGN INX12 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.45 2.50 4.05 ;
        RECT  2.00 2.45 2.50 10.55 ;
        RECT  1.80 7.45 2.50 10.55 ;
        RECT  4.45 2.45 4.95 10.55 ;
        RECT  4.45 7.45 5.20 10.55 ;
        RECT  4.45 2.45 5.35 4.95 ;
        RECT  2.00 4.45 7.70 4.95 ;
        RECT  7.20 2.45 7.70 10.55 ;
        RECT  7.20 2.45 7.90 4.05 ;
        RECT  7.20 7.45 7.90 10.55 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.30 1.15 11.00 ;
        RECT  3.15 7.30 3.85 11.00 ;
        RECT  5.85 7.30 6.55 11.00 ;
        RECT  8.55 7.30 9.25 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 4.00 ;
        RECT  3.15 2.00 3.85 4.00 ;
        RECT  5.85 2.00 6.55 4.00 ;
        RECT  8.55 2.00 9.25 4.00 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
END INX12
#MACRO INX16
#    CLASS CORE ;
#    FOREIGN INX16 0.00 0.00  ;
#    ORIGIN 0.00 0.00 ;
#    SIZE 12.60 BY 13.00 ;
#    SYMMETRY x y r90 ;
#    SITE core ;
#    PIN Q
#        DIRECTION OUTPUT ;
#        ANTENNADIFFAREA 1.0 ;
#        PORT
#        LAYER M1M ;
#        RECT  1.90 2.45 2.60 4.05 ;
#        RECT  2.10 2.45 2.60 10.55 ;
#        RECT  1.90 7.45 2.60 10.55 ;
#        RECT  4.45 2.45 5.35 4.95 ;
#        RECT  4.85 2.45 5.35 10.55 ;
#        RECT  4.60 7.45 5.35 10.55 ;
#        RECT  7.30 2.45 7.80 10.55 ;
#        RECT  7.30 2.45 8.00 4.95 ;
#        RECT  7.30 7.45 8.00 10.55 ;
#        RECT  2.10 4.45 10.50 4.95 ;
#        RECT  10.00 2.45 10.50 10.55 ;
#        RECT  10.00 2.45 10.70 4.05 ;
#        RECT  10.00 7.45 10.70 10.55 ;
#        END
#    END Q
#    PIN A
#        DIRECTION INPUT ;
#        ANTENNAGATEAREA 16.80 ;
#        PORT
#        LAYER M1M ;
#        RECT  5.85 5.40 6.75 6.30 ;
#        END
#    END A
#    PIN vdd!
#        DIRECTION INOUT ;
#        USE power ;
#        SHAPE ABUTMENT ;
#        PORT
#        LAYER M1M ;
#        RECT  0.55 7.30 1.25 11.00 ;
#        RECT  3.25 7.30 3.95 11.00 ;
#        RECT  5.95 7.30 6.65 11.00 ;
#        RECT  8.65 7.30 9.35 11.00 ;
#        RECT  11.35 7.30 12.05 11.00 ;
#        RECT  0.00 11.00 12.60 13.00 ;
#        END
#    END vdd!
#    PIN gnd!
#        DIRECTION INOUT ;
#        USE ground ;
#        SHAPE ABUTMENT ;
#        PORT
#        LAYER M1M ;
#        RECT  0.55 2.00 1.25 4.00 ;
#        RECT  3.25 2.00 3.95 4.00 ;
#        RECT  5.95 2.00 6.65 4.00 ;
#        RECT  8.65 2.00 9.35 4.00 ;
#        RECT  11.35 2.00 12.05 4.00 ;
#        RECT  0.00 0.00 12.60 2.00 ;
#        END
#    END gnd!
#END INX16
MACRO INX2
    CLASS CORE ;
    FOREIGN INX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.75 2.55 4.35 ;
        RECT  2.00 2.75 2.55 10.55 ;
        RECT  1.65 7.15 2.55 10.55 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.15 1.15 11.00 ;
        RECT  0.00 11.00 4.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 4.35 ;
        RECT  0.00 0.00 4.20 2.00 ;
        END
    END gnd!
END INX2
MACRO INX20
    CLASS CORE ;
    FOREIGN INX20 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.90 2.45 2.60 4.05 ;
        RECT  2.10 2.45 2.60 10.55 ;
        RECT  1.90 7.45 2.60 10.55 ;
        RECT  4.60 2.45 5.35 4.95 ;
        RECT  4.85 2.45 5.35 10.55 ;
        RECT  4.60 7.45 5.35 10.55 ;
        RECT  7.30 2.45 7.80 10.55 ;
        RECT  7.30 7.45 8.00 10.55 ;
        RECT  7.25 2.45 8.15 4.95 ;
        RECT  10.00 2.45 10.50 10.55 ;
        RECT  10.00 2.45 10.70 4.95 ;
        RECT  10.00 7.45 10.70 10.55 ;
        RECT  2.10 4.45 13.20 4.95 ;
        RECT  12.70 2.45 13.20 10.55 ;
        RECT  12.70 2.45 13.40 4.05 ;
        RECT  12.70 7.45 13.40 10.55 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 21.00 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.55 7.30 1.25 11.00 ;
        RECT  3.25 7.30 3.95 11.00 ;
        RECT  5.95 7.30 6.65 11.00 ;
        RECT  8.65 7.30 9.35 11.00 ;
        RECT  11.35 7.30 12.05 11.00 ;
        RECT  14.05 7.30 14.75 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.55 2.00 1.25 4.00 ;
        RECT  3.25 2.00 3.95 4.00 ;
        RECT  5.95 2.00 6.65 4.00 ;
        RECT  8.65 2.00 9.35 4.00 ;
        RECT  11.35 2.00 12.05 4.00 ;
        RECT  14.05 2.00 14.75 4.00 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
END INX20
MACRO INX3
    CLASS CORE ;
    FOREIGN INX3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.80 2.50 4.50 ;
        RECT  1.80 4.00 3.55 4.50 ;
        RECT  3.05 4.00 3.55 9.65 ;
        RECT  3.05 7.15 3.95 9.65 ;
        RECT  1.95 8.85 3.95 9.65 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.15 1.15 11.00 ;
        RECT  0.45 7.15 2.40 7.85 ;
        RECT  0.45 10.30 2.45 11.00 ;
        RECT  0.00 11.00 4.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 4.45 ;
        RECT  0.00 0.00 4.20 2.00 ;
        END
    END gnd!
END INX3
MACRO INX4
    CLASS CORE ;
    FOREIGN INX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.65 2.45 2.55 4.05 ;
        RECT  2.05 2.45 2.55 10.55 ;
        RECT  1.80 7.15 2.55 10.55 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.20 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.20 1.15 11.00 ;
        RECT  3.15 7.20 3.85 11.00 ;
        RECT  0.00 11.00 5.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 4.00 ;
        RECT  3.15 2.00 3.85 4.00 ;
        RECT  0.00 0.00 5.60 2.00 ;
        END
    END gnd!
END INX4
MACRO INX8
    CLASS CORE ;
    FOREIGN INX8 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
       DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.45 2.50 4.05 ;
        RECT  2.00 2.45 2.50 10.55 ;
        RECT  1.80 7.45 2.50 10.55 ;
        RECT  2.00 5.30 5.35 5.80 ;
        RECT  4.45 2.45 4.95 10.55 ;
        RECT  4.45 2.45 5.20 4.05 ;
        RECT  4.45 7.45 5.20 10.55 ;
        RECT  4.45 5.30 5.35 6.30 ;
        END
    END Q
#    PIN A
#        DIRECTION INPUT ;
#        ANTENNAGATEAREA 8.40 ;
#        PORT
#        LAYER M1M ;
#        RECT  0.25 5.40 1.15 6.30 ;
#        END
#    END A
#    PIN vdd!
#        DIRECTION INOUT ;
#        USE power ;
#        SHAPE ABUTMENT ;
#        PORT
#        LAYER M1M ;
#        RECT  0.45 7.70 1.15 11.00 ;
#        RECT  3.15 7.30 3.85 11.00 ;
#        RECT  5.85 7.30 6.55 11.00 ;
#        RECT  0.00 11.00 7.00 13.00 ;
#        END
#    END vdd!
#    PIN gnd!
#        DIRECTION INOUT ;
#        USE ground ;
#        SHAPE ABUTMENT ;
#        PORT
#        LAYER M1M ;
#        RECT  0.45 2.00 1.15 4.00 ;
#        RECT  3.15 2.00 3.85 4.00 ;
#        RECT  5.85 2.00 6.55 4.00 ;
#        RECT  0.00 0.00 7.00 2.00 ;
#        END
#    END gnd!
#END INX8
MACRO ITHCX12
    CLASS CORE ;
    FOREIGN ITHCX12 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.45 6.75 12.25 10.55 ;
        RECT  12.40 2.45 13.10 4.60 ;
        RECT  12.60 2.45 13.10 5.40 ;
        RECT  14.15 6.75 14.95 10.55 ;
        RECT  15.65 2.45 16.25 6.30 ;
        RECT  15.55 2.45 16.25 5.40 ;
        RECT  16.00 2.45 16.25 7.25 ;
        RECT  12.60 4.90 16.25 5.40 ;
        RECT  16.00 5.40 16.50 7.25 ;
        RECT  15.65 5.40 16.55 6.30 ;
        RECT  11.45 6.75 17.65 7.25 ;
        RECT  16.85 6.75 17.65 10.55 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.24 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.95 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.70 8.05 3.60 11.00 ;
        RECT  0.40 10.55 3.60 11.00 ;
        RECT  5.80 9.70 6.55 11.00 ;
        RECT  7.40 7.70 8.20 11.00 ;
        RECT  10.10 7.10 10.90 11.00 ;
        RECT  12.80 7.70 13.60 11.00 ;
        RECT  15.50 7.70 16.30 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.35 2.00 2.05 2.85 ;
        RECT  5.00 2.00 5.70 3.25 ;
        RECT  7.70 2.00 8.40 3.25 ;
        RECT  11.05 2.00 11.75 4.50 ;
        RECT  14.15 2.00 14.45 4.45 ;
        RECT  13.75 2.80 14.45 4.45 ;
        RECT  14.15 2.00 14.95 3.30 ;
        RECT  13.75 2.80 14.95 3.30 ;
        RECT  17.05 2.00 17.75 4.50 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.35 3.75 2.10 4.50 ;
        RECT  1.60 3.75 2.10 9.65 ;
        RECT  1.30 7.80 2.10 9.65 ;
        RECT  3.30 2.45 4.10 3.30 ;
        RECT  3.60 2.45 4.10 4.75 ;
        RECT  3.65 5.20 4.35 5.90 ;
        RECT  1.60 5.40 4.35 5.90 ;
        RECT  4.20 8.00 5.30 8.70 ;
        RECT  4.80 4.25 5.30 9.85 ;
        RECT  4.65 8.00 5.30 9.85 ;
        RECT  4.65 9.15 5.35 9.85 ;
        RECT  5.45 4.05 6.15 4.75 ;
        RECT  3.60 4.25 6.15 4.75 ;
        RECT  5.75 6.75 6.55 7.85 ;
        RECT  6.30 2.45 7.10 3.40 ;
        RECT  6.60 2.45 7.10 4.95 ;
        RECT  7.20 4.45 7.70 7.25 ;
        RECT  5.75 6.75 7.70 7.25 ;
        RECT  6.60 4.45 9.10 4.95 ;
        RECT  8.40 4.45 9.10 5.25 ;
        RECT  9.05 5.85 9.55 10.55 ;
        RECT  8.75 7.05 9.55 10.55 ;
        RECT  9.55 3.55 10.30 4.30 ;
        RECT  9.80 3.55 10.30 6.35 ;
        RECT  9.80 5.65 11.20 6.35 ;
        RECT  9.05 5.85 11.20 6.35 ;
    END
END ITHCX12
MACRO ITHCX16
    CLASS CORE ;
    FOREIGN ITHCX16 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  14.35 6.80 15.15 10.55 ;
        RECT  15.75 2.45 16.45 4.60 ;
        RECT  15.95 2.45 16.45 5.40 ;
        RECT  17.05 6.80 17.85 10.55 ;
        RECT  18.45 2.45 19.20 5.40 ;
        RECT  19.90 6.80 20.70 10.55 ;
        RECT  21.15 2.45 21.90 5.40 ;
        RECT  21.25 2.45 21.90 6.30 ;
        RECT  21.25 5.40 22.15 6.30 ;
        RECT  21.65 2.45 21.90 7.30 ;
        RECT  15.95 4.90 21.90 5.40 ;
        RECT  21.65 5.40 22.15 7.30 ;
        RECT  14.35 6.80 23.40 7.30 ;
        RECT  22.60 6.80 23.40 10.55 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.85 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.50 2.55 7.60 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.33 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.75 8.30 2.55 11.00 ;
        RECT  3.45 7.20 3.95 11.00 ;
        RECT  3.45 7.20 4.45 9.05 ;
        RECT  7.65 7.40 8.40 11.00 ;
        RECT  10.30 7.70 11.10 11.00 ;
        RECT  13.00 7.75 13.80 11.00 ;
        RECT  15.70 7.75 16.50 11.00 ;
        RECT  18.45 7.75 19.30 11.00 ;
        RECT  21.25 7.75 22.05 11.00 ;
        RECT  0.00 11.00 23.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.75 2.00 2.55 3.15 ;
        RECT  5.35 2.00 6.05 4.40 ;
        RECT  5.35 2.00 7.25 2.25 ;
        RECT  9.25 2.00 9.95 4.00 ;
        RECT  11.00 2.00 13.55 2.10 ;
        RECT  14.40 2.00 15.10 4.50 ;
        RECT  17.10 2.00 17.80 4.45 ;
        RECT  19.80 2.00 20.50 4.45 ;
        RECT  22.65 2.00 23.35 4.50 ;
        RECT  0.00 0.00 23.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.30 4.85 5.45 5.45 ;
        RECT  0.70 5.90 4.10 6.05 ;
        RECT  0.70 5.55 1.20 10.55 ;
        RECT  0.45 8.35 1.20 10.55 ;
        RECT  1.80 3.80 2.30 6.05 ;
        RECT  1.80 3.80 2.50 4.50 ;
        RECT  3.35 5.55 3.85 6.70 ;
        RECT  0.70 5.55 3.85 6.05 ;
        RECT  3.35 5.90 4.10 6.70 ;
        RECT  3.70 2.90 4.90 3.60 ;
        RECT  4.40 2.90 4.90 5.45 ;
        RECT  4.95 4.75 5.05 10.25 ;
        RECT  4.30 4.75 5.05 5.45 ;
        RECT  4.95 4.85 5.45 10.25 ;
        RECT  4.40 9.50 5.45 10.25 ;
        RECT  4.40 9.75 6.65 10.25 ;
        RECT  5.90 9.75 6.65 10.55 ;
        RECT  6.70 2.80 7.20 8.85 ;
        RECT  6.05 7.25 7.20 8.85 ;
        RECT  6.70 2.80 7.40 4.95 ;
        RECT  7.90 2.55 8.60 3.30 ;
        RECT  6.70 2.80 8.60 3.30 ;
        RECT  8.95 6.75 9.75 10.55 ;
        RECT  6.70 4.45 12.85 4.95 ;
        RECT  11.75 3.30 12.45 4.00 ;
        RECT  12.00 5.85 12.45 10.55 ;
        RECT  11.65 6.75 12.45 10.55 ;
        RECT  12.00 5.85 12.50 7.25 ;
        RECT  8.95 6.75 12.50 7.25 ;
        RECT  12.15 4.45 12.85 5.15 ;
        RECT  11.75 3.50 13.95 4.00 ;
        RECT  13.45 3.50 13.95 6.35 ;
        RECT  13.45 5.65 14.20 6.35 ;
        RECT  12.00 5.85 14.20 6.35 ;
    END
END ITHCX16
MACRO ITHCX20
    CLASS CORE ;
    FOREIGN ITHCX20 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 25.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  14.35 6.80 15.15 10.55 ;
        RECT  15.75 2.45 16.45 4.60 ;
        RECT  15.95 2.45 16.45 5.40 ;
        RECT  17.05 6.80 17.85 10.55 ;
        RECT  18.45 2.45 19.20 5.40 ;
        RECT  19.75 6.80 20.55 10.55 ;
        RECT  21.15 2.45 21.90 5.40 ;
        RECT  21.25 2.45 21.90 6.30 ;
        RECT  21.25 5.40 22.15 6.30 ;
        RECT  21.65 2.45 21.90 7.30 ;
        RECT  15.95 4.90 21.90 5.40 ;
        RECT  21.65 5.40 22.15 7.30 ;
        RECT  14.35 6.80 23.25 7.30 ;
        RECT  22.45 6.80 23.25 10.55 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.85 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.50 2.55 7.60 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.33 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.75 8.30 2.55 11.00 ;
        RECT  3.45 7.20 3.95 11.00 ;
        RECT  3.45 7.20 4.45 9.05 ;
        RECT  7.65 7.40 8.40 11.00 ;
        RECT  10.30 7.70 11.10 11.00 ;
        RECT  13.00 7.75 13.80 11.00 ;
        RECT  15.70 7.75 16.50 11.00 ;
        RECT  18.45 7.75 19.15 11.00 ;
        RECT  21.10 7.75 21.90 11.00 ;
        RECT  23.95 6.90 24.75 11.00 ;
        RECT  0.00 11.00 25.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.60 2.00 2.40 3.15 ;
        RECT  5.35 2.00 6.05 4.40 ;
        RECT  5.35 2.00 7.25 2.25 ;
        RECT  9.25 2.00 9.95 4.00 ;
        RECT  11.00 2.00 13.55 2.10 ;
        RECT  14.40 2.00 15.10 4.50 ;
        RECT  17.10 2.00 17.80 4.45 ;
        RECT  19.80 2.00 20.50 4.45 ;
        RECT  22.50 2.00 23.20 4.55 ;
        RECT  24.05 2.00 24.75 4.50 ;
        RECT  0.00 0.00 25.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.30 4.85 5.45 5.45 ;
        RECT  0.70 5.90 4.10 6.05 ;
        RECT  0.70 5.55 1.20 10.55 ;
        RECT  0.45 8.35 1.20 10.55 ;
        RECT  1.60 3.80 2.10 6.05 ;
        RECT  1.60 3.80 2.30 4.50 ;
        RECT  3.35 5.55 3.85 6.70 ;
        RECT  0.70 5.55 3.85 6.05 ;
        RECT  3.35 5.90 4.10 6.70 ;
        RECT  3.70 2.90 4.90 3.60 ;
        RECT  4.40 2.90 4.90 5.45 ;
        RECT  4.95 4.75 5.05 10.25 ;
        RECT  4.30 4.75 5.05 5.45 ;
        RECT  4.95 4.85 5.45 10.25 ;
        RECT  4.40 9.50 5.45 10.25 ;
        RECT  4.40 9.75 6.65 10.25 ;
        RECT  5.90 9.75 6.65 10.55 ;
        RECT  6.70 2.80 7.20 8.85 ;
        RECT  6.05 7.25 7.20 8.85 ;
        RECT  6.70 2.80 7.40 4.95 ;
        RECT  7.90 2.55 8.60 3.30 ;
        RECT  6.70 2.80 8.60 3.30 ;
        RECT  8.95 6.75 9.75 10.55 ;
        RECT  6.70 4.45 12.85 4.95 ;
        RECT  11.75 3.30 12.45 4.00 ;
        RECT  12.00 5.85 12.45 10.55 ;
        RECT  11.65 6.75 12.45 10.55 ;
        RECT  12.00 5.85 12.50 7.25 ;
        RECT  8.95 6.75 12.50 7.25 ;
        RECT  12.15 4.45 12.85 5.15 ;
        RECT  11.75 3.50 13.95 4.00 ;
        RECT  13.45 3.50 13.95 6.35 ;
        RECT  13.45 5.65 14.20 6.35 ;
        RECT  12.00 5.85 14.20 6.35 ;
    END
END ITHCX20
MACRO ITHCX3
    CLASS CORE ;
    FOREIGN ITHCX3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.30 6.75 10.80 10.55 ;
        RECT  10.00 7.95 10.80 10.55 ;
        RECT  11.40 2.45 12.10 4.60 ;
        RECT  11.65 2.45 12.10 7.25 ;
        RECT  11.60 2.45 12.10 6.30 ;
        RECT  11.65 5.40 12.15 7.25 ;
        RECT  10.30 6.75 12.15 7.25 ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.58 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.55 7.60 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.67 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 8.05 2.70 11.00 ;
        RECT  0.40 10.85 2.70 11.00 ;
        RECT  5.95 8.90 6.75 11.00 ;
        RECT  4.85 9.70 6.75 11.00 ;
        RECT  8.65 9.05 9.45 11.00 ;
        RECT  11.35 7.95 12.15 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.55 2.00 3.25 2.25 ;
        RECT  4.15 2.00 4.95 4.25 ;
        RECT  6.85 2.00 7.65 4.40 ;
        RECT  10.05 2.00 10.75 4.50 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.90 2.65 2.10 3.15 ;
        RECT  0.25 5.65 0.75 9.75 ;
        RECT  0.25 8.75 1.20 9.75 ;
        RECT  0.90 2.45 1.60 3.15 ;
        RECT  1.60 2.65 2.10 6.15 ;
        RECT  2.55 3.20 3.40 3.90 ;
        RECT  0.25 5.65 3.65 6.15 ;
        RECT  2.90 3.20 3.40 5.20 ;
        RECT  2.90 4.25 3.60 5.20 ;
        RECT  2.95 5.65 3.65 6.35 ;
        RECT  2.90 4.70 4.60 5.20 ;
        RECT  4.10 4.70 4.15 9.85 ;
        RECT  3.35 7.75 4.15 9.85 ;
        RECT  3.35 9.15 4.40 9.85 ;
        RECT  4.10 4.70 4.60 8.25 ;
        RECT  3.35 7.75 4.60 8.25 ;
        RECT  5.50 3.50 6.35 4.40 ;
        RECT  5.85 3.50 6.35 7.80 ;
        RECT  5.05 7.10 6.35 7.80 ;
        RECT  7.30 5.45 8.00 6.15 ;
        RECT  5.85 5.65 8.00 6.15 ;
        RECT  7.60 7.30 8.10 10.55 ;
        RECT  7.30 8.95 8.10 10.55 ;
        RECT  8.50 3.70 9.30 4.45 ;
        RECT  8.80 3.70 9.30 7.80 ;
        RECT  7.60 7.30 9.30 7.80 ;
        RECT  8.80 6.80 9.85 7.50 ;
        RECT  7.60 7.30 9.85 7.50 ;
    END
END ITHCX3
MACRO ITHCX4
    CLASS CORE ;
    FOREIGN ITHCX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.30 6.75 10.80 10.55 ;
        RECT  10.00 7.95 10.80 10.55 ;
        RECT  11.25 2.45 11.95 4.60 ;
        RECT  11.75 2.45 11.95 7.25 ;
        RECT  11.45 2.45 11.95 6.30 ;
        RECT  11.75 5.40 12.25 7.25 ;
        RECT  10.30 6.75 12.25 7.25 ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.58 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.55 7.60 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.67 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.05 2.70 11.00 ;
        RECT  5.85 8.90 6.70 11.00 ;
        RECT  4.85 9.70 6.70 11.00 ;
        RECT  8.65 8.95 9.45 11.00 ;
        RECT  11.35 7.95 12.15 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.75 2.00 3.45 2.60 ;
        RECT  4.15 2.00 4.95 4.25 ;
        RECT  6.85 2.00 7.65 4.40 ;
        RECT  9.90 2.00 10.60 4.50 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.25 5.75 0.75 9.85 ;
        RECT  0.25 9.15 1.15 9.85 ;
        RECT  0.95 2.80 2.10 3.50 ;
        RECT  1.60 2.80 2.10 6.25 ;
        RECT  2.65 3.55 3.50 4.35 ;
        RECT  0.25 5.75 3.65 6.25 ;
        RECT  2.95 3.55 3.50 5.20 ;
        RECT  2.95 5.65 3.65 6.35 ;
        RECT  3.35 7.95 4.20 8.65 ;
        RECT  2.95 4.70 4.90 5.20 ;
        RECT  4.10 4.70 4.20 9.85 ;
        RECT  3.70 7.95 4.20 9.85 ;
        RECT  3.70 9.15 4.40 9.85 ;
        RECT  4.10 4.70 4.60 8.45 ;
        RECT  3.35 7.95 4.60 8.45 ;
        RECT  4.10 4.70 4.90 5.40 ;
        RECT  5.50 3.50 6.30 4.40 ;
        RECT  5.80 3.50 6.30 7.80 ;
        RECT  5.05 7.10 6.30 7.80 ;
        RECT  7.60 7.00 8.10 10.55 ;
        RECT  7.30 8.95 8.10 10.55 ;
        RECT  7.45 5.45 8.15 6.15 ;
        RECT  5.80 5.65 8.15 6.15 ;
        RECT  8.40 3.70 9.10 4.45 ;
        RECT  8.60 3.70 9.10 7.50 ;
        RECT  8.60 6.80 9.85 7.50 ;
        RECT  7.60 7.00 9.85 7.50 ;
    END
END ITHCX4
MACRO ITHCX8
    CLASS CORE ;
    FOREIGN ITHCX8 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.45 6.75 12.25 10.55 ;
        RECT  12.40 2.45 13.10 4.60 ;
        RECT  12.60 2.45 13.10 6.30 ;
        RECT  13.20 5.40 13.70 7.25 ;
        RECT  12.60 5.40 13.75 6.30 ;
        RECT  11.45 6.75 14.95 7.25 ;
        RECT  14.15 6.75 14.95 10.55 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.24 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.95 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.70 8.05 3.60 11.00 ;
        RECT  0.40 10.55 3.60 11.00 ;
        RECT  5.80 9.70 6.55 11.00 ;
        RECT  7.40 7.70 8.20 11.00 ;
        RECT  10.10 7.10 10.90 11.00 ;
        RECT  12.80 7.70 13.60 11.00 ;
        RECT  15.50 7.70 16.30 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.35 2.00 2.05 2.85 ;
        RECT  5.00 2.00 5.70 3.25 ;
        RECT  7.70 2.00 8.40 3.25 ;
        RECT  11.05 2.00 11.75 4.50 ;
        RECT  14.10 2.00 14.85 4.45 ;
        RECT  13.75 3.40 14.85 4.45 ;
        RECT  15.65 2.00 16.35 4.50 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.35 3.75 2.10 4.50 ;
        RECT  1.60 3.75 2.10 9.65 ;
        RECT  1.30 7.80 2.10 9.65 ;
        RECT  3.30 2.45 4.10 3.30 ;
        RECT  3.60 2.45 4.10 4.75 ;
        RECT  3.65 5.20 4.35 5.90 ;
        RECT  1.60 5.40 4.35 5.90 ;
        RECT  4.20 8.00 5.30 8.70 ;
        RECT  4.80 4.25 5.30 9.85 ;
        RECT  4.65 8.00 5.30 9.85 ;
        RECT  4.65 9.15 5.35 9.85 ;
        RECT  5.45 4.05 6.15 4.75 ;
        RECT  3.60 4.25 6.15 4.75 ;
        RECT  5.75 6.75 6.55 7.85 ;
        RECT  6.30 2.45 7.10 3.40 ;
        RECT  6.60 2.45 7.10 4.95 ;
        RECT  7.20 4.45 7.70 7.25 ;
        RECT  5.75 6.75 7.70 7.25 ;
        RECT  6.60 4.45 9.10 4.95 ;
        RECT  8.40 4.45 9.10 5.25 ;
        RECT  9.05 5.85 9.55 10.55 ;
        RECT  8.75 7.05 9.55 10.55 ;
        RECT  9.55 3.55 10.30 4.30 ;
        RECT  9.80 3.55 10.30 6.35 ;
        RECT  9.80 5.65 11.20 6.35 ;
        RECT  9.05 5.85 11.20 6.35 ;
    END
END ITHCX8
MACRO ITHX1
    CLASS CORE ;
    FOREIGN ITHX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.30 2.70 5.35 4.45 ;
        RECT  4.85 2.70 5.35 10.55 ;
        RECT  4.30 7.70 5.35 10.55 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 9.30 1.15 10.20 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 3.10 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.95 7.70 2.65 11.00 ;
        RECT  0.00 11.00 5.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.95 2.00 2.65 4.45 ;
        RECT  0.00 0.00 5.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.75 0.95 8.85 ;
        RECT  0.45 3.75 1.15 4.45 ;
        RECT  0.45 6.75 1.15 8.85 ;
        RECT  3.65 6.10 4.35 7.25 ;
        RECT  0.45 6.75 4.35 7.25 ;
    END
END ITHX1
MACRO ITHX12
    CLASS CORE ;
    FOREIGN ITHX12 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.65 8.00 9.55 8.90 ;
        RECT  8.80 2.45 9.55 4.05 ;
        RECT  9.00 2.45 9.55 10.55 ;
        RECT  8.80 7.70 9.55 10.55 ;
        RECT  11.50 6.50 12.00 10.55 ;
        RECT  11.50 2.45 12.20 4.90 ;
        RECT  11.50 7.70 12.20 10.55 ;
        RECT  9.00 6.50 14.70 7.00 ;
        RECT  14.20 2.45 14.70 4.90 ;
        RECT  9.00 4.40 14.70 4.90 ;
        RECT  14.20 6.50 14.70 10.55 ;
        RECT  14.20 2.45 14.90 4.05 ;
        RECT  14.20 7.70 14.90 10.55 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.65 9.25 1.35 11.00 ;
        RECT  4.60 9.95 5.30 11.00 ;
        RECT  7.45 7.70 8.15 11.00 ;
        RECT  10.15 7.55 10.85 11.00 ;
        RECT  12.85 7.55 13.55 11.00 ;
        RECT  15.55 7.70 16.25 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.60 ;
        RECT  7.45 2.00 8.15 4.00 ;
        RECT  10.15 2.00 10.85 3.95 ;
        RECT  12.85 2.00 13.55 3.95 ;
        RECT  15.55 2.00 16.25 4.00 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.60 6.05 2.35 6.75 ;
        RECT  2.80 6.85 3.95 7.35 ;
        RECT  0.95 3.25 2.10 3.95 ;
        RECT  1.85 3.25 2.10 10.45 ;
        RECT  1.60 3.25 2.10 6.75 ;
        RECT  1.85 6.05 2.35 10.45 ;
        RECT  1.85 9.75 2.70 10.45 ;
        RECT  2.55 3.45 3.30 4.15 ;
        RECT  3.25 3.45 3.30 9.50 ;
        RECT  2.80 3.45 3.30 7.35 ;
        RECT  3.25 6.85 3.95 9.50 ;
        RECT  4.10 2.55 4.80 4.95 ;
        RECT  4.80 4.45 5.30 8.55 ;
        RECT  4.60 6.85 5.30 8.55 ;
        RECT  3.25 9.00 6.80 9.50 ;
        RECT  6.10 2.45 6.80 4.95 ;
        RECT  6.30 6.75 6.80 10.55 ;
        RECT  6.10 7.70 6.80 10.55 ;
        RECT  4.10 4.45 8.50 4.95 ;
        RECT  7.80 4.45 8.50 5.15 ;
        RECT  7.85 6.50 8.55 7.25 ;
        RECT  6.30 6.75 8.55 7.25 ;
        RECT  10.00 5.35 10.70 6.05 ;
        RECT  10.00 5.55 16.60 6.05 ;
        RECT  16.10 4.45 16.60 7.25 ;
        RECT  16.10 6.75 17.55 7.25 ;
        RECT  17.05 3.35 17.55 4.95 ;
        RECT  16.10 4.45 17.55 4.95 ;
        RECT  17.05 6.75 17.55 9.40 ;
        RECT  17.05 3.35 17.75 4.05 ;
        RECT  17.05 7.70 17.75 9.40 ;
    END
END ITHX12
MACRO ITHX16
    CLASS CORE ;
    FOREIGN ITHX16 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.65 2.80 9.60 3.70 ;
        RECT  8.90 2.45 9.60 4.05 ;
        RECT  9.30 2.45 9.60 10.55 ;
        RECT  9.10 2.45 9.60 4.90 ;
        RECT  9.30 4.40 9.80 10.55 ;
        RECT  9.00 7.70 9.80 10.55 ;
        RECT  11.60 2.45 12.30 4.90 ;
        RECT  11.70 6.50 12.40 10.55 ;
        RECT  14.30 2.45 15.00 4.90 ;
        RECT  14.40 6.50 15.10 10.55 ;
        RECT  9.30 6.50 17.60 7.00 ;
        RECT  17.00 2.45 17.50 4.90 ;
        RECT  9.10 4.40 17.50 4.90 ;
        RECT  17.10 6.50 17.60 10.55 ;
        RECT  17.00 2.45 17.70 4.05 ;
        RECT  17.10 7.70 17.80 10.55 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.65 9.25 1.35 11.00 ;
        RECT  4.35 9.95 5.05 11.00 ;
        RECT  7.65 7.70 8.35 11.00 ;
        RECT  10.35 7.55 11.05 11.00 ;
        RECT  13.05 7.55 13.75 11.00 ;
        RECT  15.75 7.55 16.45 11.00 ;
        RECT  18.45 7.70 19.15 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.60 ;
        RECT  7.40 2.00 8.10 4.00 ;
        RECT  10.25 2.00 10.95 3.95 ;
        RECT  12.95 2.00 13.65 3.95 ;
        RECT  15.65 2.00 16.35 3.95 ;
        RECT  18.35 2.00 19.05 4.00 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.60 6.05 2.35 6.75 ;
        RECT  2.80 6.85 3.70 7.35 ;
        RECT  0.95 3.25 2.10 3.95 ;
        RECT  1.85 3.25 2.10 10.55 ;
        RECT  1.60 3.25 2.10 6.75 ;
        RECT  1.85 6.05 2.35 10.55 ;
        RECT  1.85 9.85 2.70 10.55 ;
        RECT  2.55 3.45 3.30 4.15 ;
        RECT  3.00 3.45 3.30 9.50 ;
        RECT  2.80 3.45 3.30 7.35 ;
        RECT  3.00 6.85 3.70 9.50 ;
        RECT  4.55 2.55 4.80 8.55 ;
        RECT  4.10 2.55 4.80 4.95 ;
        RECT  4.55 4.45 5.05 8.55 ;
        RECT  4.35 6.85 5.05 8.55 ;
        RECT  3.00 9.00 6.75 9.50 ;
        RECT  6.05 2.45 6.75 4.95 ;
        RECT  6.25 6.75 6.75 10.55 ;
        RECT  6.05 8.05 6.75 10.55 ;
        RECT  4.10 4.45 8.65 4.95 ;
        RECT  7.95 4.45 8.65 5.15 ;
        RECT  8.15 6.50 8.85 7.25 ;
        RECT  6.25 6.75 8.85 7.25 ;
        RECT  10.25 5.35 10.95 6.05 ;
        RECT  10.25 5.55 19.40 6.05 ;
        RECT  18.90 4.45 19.40 7.25 ;
        RECT  18.90 6.75 20.35 7.25 ;
        RECT  19.85 3.35 20.35 4.95 ;
        RECT  18.90 4.45 20.35 4.95 ;
        RECT  19.85 6.75 20.35 9.40 ;
        RECT  19.85 3.35 20.55 4.05 ;
        RECT  19.85 7.70 20.55 9.40 ;
    END
END ITHX16
MACRO ITHX2
    CLASS CORE ;
    FOREIGN ITHX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.80 2.45 9.30 10.55 ;
        RECT  8.60 7.80 9.30 10.55 ;
        RECT  8.65 2.45 9.55 4.05 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.45 1.15 11.00 ;
        RECT  4.40 10.25 5.10 11.00 ;
        RECT  7.25 7.80 7.95 11.00 ;
        RECT  11.45 7.15 12.15 11.00 ;
        RECT  10.25 10.10 12.15 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.75 ;
        RECT  7.35 2.00 8.05 4.00 ;
        RECT  10.40 2.00 11.10 3.15 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.80 5.40 3.80 5.90 ;
        RECT  0.95 3.40 2.10 4.10 ;
        RECT  1.80 3.40 2.10 9.15 ;
        RECT  1.60 3.40 2.10 7.05 ;
        RECT  1.80 6.35 2.50 9.15 ;
        RECT  2.60 3.60 3.30 4.30 ;
        RECT  1.60 6.35 2.85 7.05 ;
        RECT  2.80 3.60 3.30 5.90 ;
        RECT  3.30 5.40 3.80 9.80 ;
        RECT  3.30 7.15 4.00 9.80 ;
        RECT  4.65 2.70 4.85 8.85 ;
        RECT  4.15 2.70 4.85 4.95 ;
        RECT  4.65 4.45 5.15 8.85 ;
        RECT  4.65 7.15 5.35 8.85 ;
        RECT  3.30 9.30 6.45 9.80 ;
        RECT  5.95 6.85 6.45 10.55 ;
        RECT  5.75 9.30 6.45 10.55 ;
        RECT  5.85 3.35 6.55 4.95 ;
        RECT  4.15 4.45 8.35 4.95 ;
        RECT  7.65 4.45 8.35 5.15 ;
        RECT  7.65 6.65 8.35 7.35 ;
        RECT  5.95 6.85 8.35 7.35 ;
        RECT  9.75 5.85 10.80 6.55 ;
        RECT  10.30 3.80 10.80 8.85 ;
        RECT  10.10 5.85 10.80 8.85 ;
        RECT  10.30 3.80 11.10 4.50 ;
    END
END ITHX2
MACRO ITHX20
    CLASS CORE ;
    FOREIGN ITHX20 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  9.00 2.45 9.75 4.05 ;
        RECT  9.55 2.45 9.75 10.55 ;
        RECT  9.25 2.45 9.75 4.90 ;
        RECT  9.55 4.40 10.05 10.55 ;
        RECT  9.15 7.75 10.05 10.55 ;
        RECT  11.70 2.45 12.40 4.90 ;
        RECT  11.85 6.50 12.55 10.55 ;
        RECT  14.40 2.45 15.10 4.90 ;
        RECT  14.55 6.50 15.25 10.55 ;
        RECT  17.05 6.50 17.95 7.60 ;
        RECT  17.10 2.45 17.80 4.90 ;
        RECT  17.25 6.50 17.95 10.55 ;
        RECT  9.55 6.50 20.65 7.00 ;
        RECT  19.80 2.45 20.50 4.90 ;
        RECT  9.25 4.40 20.50 4.90 ;
        RECT  19.95 6.50 20.65 10.55 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  22.65 5.40 23.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 9.45 1.15 11.00 ;
        RECT  3.35 9.95 4.05 11.00 ;
        RECT  7.75 7.75 8.45 11.00 ;
        RECT  10.50 7.45 11.20 11.00 ;
        RECT  13.20 7.45 13.90 11.00 ;
        RECT  15.90 7.45 16.60 11.00 ;
        RECT  18.60 7.45 19.30 11.00 ;
        RECT  21.30 7.70 22.00 11.00 ;
        RECT  0.00 11.00 23.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.60 ;
        RECT  7.65 2.00 8.35 4.00 ;
        RECT  10.35 2.00 11.05 3.95 ;
        RECT  13.05 2.00 13.75 3.95 ;
        RECT  15.75 2.00 16.45 3.95 ;
        RECT  18.45 2.00 19.15 3.95 ;
        RECT  21.15 2.00 21.85 4.00 ;
        RECT  0.00 0.00 23.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.15 4.45 2.10 4.95 ;
        RECT  0.95 3.25 1.65 3.95 ;
        RECT  1.60 3.25 1.65 10.55 ;
        RECT  1.15 3.25 1.65 4.95 ;
        RECT  1.60 4.45 2.10 10.55 ;
        RECT  1.60 5.60 2.35 6.30 ;
        RECT  1.60 9.85 2.50 10.55 ;
        RECT  2.50 3.45 3.30 4.15 ;
        RECT  2.55 6.85 3.30 8.55 ;
        RECT  2.80 3.45 3.30 9.50 ;
        RECT  4.05 2.50 4.60 8.55 ;
        RECT  3.90 6.85 4.60 8.55 ;
        RECT  2.80 9.00 5.20 9.50 ;
        RECT  4.05 2.50 4.75 4.95 ;
        RECT  4.70 9.00 5.20 10.55 ;
        RECT  5.85 2.45 7.00 3.15 ;
        RECT  5.45 7.90 7.00 8.60 ;
        RECT  6.30 7.90 7.00 10.55 ;
        RECT  6.30 2.45 7.00 4.95 ;
        RECT  6.50 6.80 7.00 10.55 ;
        RECT  4.70 9.85 7.00 10.55 ;
        RECT  4.05 4.45 8.75 4.95 ;
        RECT  8.05 4.45 8.75 5.25 ;
        RECT  8.35 6.60 9.10 7.30 ;
        RECT  6.50 6.80 9.10 7.30 ;
        RECT  10.50 5.35 11.20 6.05 ;
        RECT  10.50 5.55 22.20 6.05 ;
        RECT  21.70 4.45 22.20 7.25 ;
        RECT  21.70 6.75 23.15 7.25 ;
        RECT  22.65 3.35 23.15 4.95 ;
        RECT  21.70 4.45 23.15 4.95 ;
        RECT  22.65 6.75 23.15 9.40 ;
        RECT  22.65 3.35 23.35 4.05 ;
        RECT  22.65 7.70 23.35 9.40 ;
    END
END ITHX20
MACRO ITHX3
    CLASS CORE ;
    FOREIGN ITHX3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.80 2.80 9.30 10.20 ;
        RECT  8.60 7.60 9.35 10.20 ;
        RECT  8.65 2.80 9.55 3.70 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  10.05 4.10 11.20 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.45 1.15 11.00 ;
        RECT  4.40 10.25 5.10 11.00 ;
        RECT  7.25 7.70 7.95 11.00 ;
        RECT  7.10 9.75 7.95 11.00 ;
        RECT  9.95 7.40 10.65 11.00 ;
        RECT  9.95 10.10 12.15 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.75 ;
        RECT  7.35 2.00 8.05 3.55 ;
        RECT  10.05 2.00 10.75 3.30 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.80 5.30 3.80 5.80 ;
        RECT  0.95 3.40 2.10 4.10 ;
        RECT  1.80 3.40 2.10 9.15 ;
        RECT  1.60 3.40 2.10 7.05 ;
        RECT  1.80 6.35 2.50 9.15 ;
        RECT  2.60 3.60 3.30 4.30 ;
        RECT  1.60 6.35 2.85 7.05 ;
        RECT  2.80 3.60 3.30 5.80 ;
        RECT  3.30 5.30 3.80 9.80 ;
        RECT  3.30 7.15 4.00 9.80 ;
        RECT  4.65 2.70 4.85 8.85 ;
        RECT  4.15 2.70 4.85 4.70 ;
        RECT  4.65 4.20 5.15 8.85 ;
        RECT  4.65 7.15 5.35 8.85 ;
        RECT  3.30 9.30 6.45 9.80 ;
        RECT  5.95 6.45 6.45 10.55 ;
        RECT  5.75 9.30 6.45 10.55 ;
        RECT  5.85 3.10 6.55 4.70 ;
        RECT  4.15 4.20 8.35 4.70 ;
        RECT  7.65 4.20 8.35 4.90 ;
        RECT  7.65 6.25 8.35 6.95 ;
        RECT  5.95 6.45 8.35 6.95 ;
        RECT  9.75 5.45 10.45 6.15 ;
        RECT  11.45 2.60 12.15 3.30 ;
        RECT  9.75 5.45 12.15 5.95 ;
        RECT  11.65 2.60 12.15 9.00 ;
        RECT  11.45 7.40 12.15 9.00 ;
    END
END ITHX3
MACRO ITHX4
    CLASS CORE ;
    FOREIGN ITHX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.60 2.45 9.30 4.05 ;
        RECT  8.80 2.45 9.30 10.55 ;
        RECT  8.60 7.70 9.30 10.55 ;
        RECT  8.60 7.70 9.55 8.90 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  11.45 9.30 12.35 10.20 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.45 1.15 11.00 ;
        RECT  4.40 10.25 5.10 11.00 ;
        RECT  7.25 7.70 7.95 11.00 ;
        RECT  10.10 7.25 10.80 11.00 ;
        RECT  9.95 9.75 10.80 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.75 ;
        RECT  7.25 2.00 7.95 4.00 ;
        RECT  9.95 2.00 10.65 4.00 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.45 4.55 2.10 5.05 ;
        RECT  0.95 3.40 1.95 4.10 ;
        RECT  1.80 3.40 1.95 9.15 ;
        RECT  1.45 3.40 1.95 5.05 ;
        RECT  1.80 4.55 2.10 9.15 ;
        RECT  1.60 4.55 2.10 7.05 ;
        RECT  1.80 6.35 2.50 9.15 ;
        RECT  2.50 3.60 3.25 4.30 ;
        RECT  1.60 6.35 2.85 7.05 ;
        RECT  2.75 3.60 3.25 5.90 ;
        RECT  2.75 5.40 3.80 5.90 ;
        RECT  3.30 5.40 3.80 9.80 ;
        RECT  3.30 7.15 4.00 9.80 ;
        RECT  4.65 2.70 4.75 8.85 ;
        RECT  4.05 2.70 4.75 4.95 ;
        RECT  4.65 4.45 5.20 8.85 ;
        RECT  4.65 7.15 5.35 8.85 ;
        RECT  3.30 9.30 6.45 9.80 ;
        RECT  5.75 3.35 6.45 4.95 ;
        RECT  5.95 6.75 6.45 10.55 ;
        RECT  5.75 9.30 6.45 10.55 ;
        RECT  4.05 4.45 8.35 4.95 ;
        RECT  7.65 4.45 8.35 5.15 ;
        RECT  7.65 6.55 8.35 7.25 ;
        RECT  5.95 6.75 8.35 7.25 ;
        RECT  9.75 5.25 11.95 5.95 ;
        RECT  11.45 3.35 11.95 8.85 ;
        RECT  11.45 3.35 12.15 4.05 ;
        RECT  11.45 7.25 12.15 8.85 ;
    END
END ITHX4
MACRO ITHX8
    CLASS CORE ;
    FOREIGN ITHX8 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.65 2.45 9.55 4.05 ;
        RECT  9.05 2.45 9.55 10.55 ;
        RECT  8.80 7.70 9.55 10.55 ;
        RECT  9.05 6.55 11.90 7.05 ;
        RECT  11.40 2.45 11.90 4.90 ;
        RECT  9.05 4.40 11.90 4.90 ;
        RECT  11.40 6.55 11.90 10.55 ;
        RECT  11.40 2.45 12.10 4.05 ;
        RECT  11.40 7.70 12.20 10.55 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.65 9.25 1.35 11.00 ;
        RECT  4.60 9.95 5.30 11.00 ;
        RECT  7.45 7.70 8.15 11.00 ;
        RECT  10.15 7.55 10.85 11.00 ;
        RECT  12.85 7.70 13.55 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.60 ;
        RECT  7.35 2.00 8.05 4.00 ;
        RECT  10.05 2.00 10.75 3.95 ;
        RECT  12.75 2.00 13.45 4.00 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.60 6.05 2.35 6.75 ;
        RECT  2.80 6.85 3.95 7.35 ;
        RECT  0.95 3.25 2.10 3.95 ;
        RECT  1.85 3.25 2.10 10.45 ;
        RECT  1.60 3.25 2.10 6.75 ;
        RECT  1.85 6.05 2.35 10.45 ;
        RECT  1.85 9.75 2.70 10.45 ;
        RECT  2.55 3.45 3.30 4.15 ;
        RECT  3.25 3.45 3.30 9.50 ;
        RECT  2.80 3.45 3.30 7.35 ;
        RECT  3.25 6.85 3.95 9.50 ;
        RECT  4.10 2.55 4.80 4.95 ;
        RECT  4.80 4.45 5.30 8.55 ;
        RECT  4.60 6.85 5.30 8.55 ;
        RECT  3.25 9.00 6.80 9.50 ;
        RECT  6.00 2.45 6.70 4.95 ;
        RECT  6.30 6.75 6.80 10.55 ;
        RECT  6.10 7.70 6.80 10.55 ;
        RECT  4.10 4.45 8.40 4.95 ;
        RECT  7.70 4.45 8.40 5.15 ;
        RECT  7.90 6.50 8.60 7.25 ;
        RECT  6.30 6.75 8.60 7.25 ;
        RECT  10.00 5.35 10.70 6.05 ;
        RECT  10.00 5.55 13.80 6.05 ;
        RECT  13.30 4.45 13.80 7.25 ;
        RECT  13.30 6.75 14.75 7.25 ;
        RECT  14.25 3.35 14.75 4.95 ;
        RECT  13.30 4.45 14.75 4.95 ;
        RECT  14.25 6.75 14.75 9.40 ;
        RECT  14.25 3.35 14.95 4.05 ;
        RECT  14.25 7.70 14.95 9.40 ;
    END
END ITHX8
MACRO ITLCX12
    CLASS CORE ;
    FOREIGN ITLCX12 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.45 6.75 12.25 10.55 ;
        RECT  12.35 2.45 13.05 4.50 ;
        RECT  12.85 2.45 13.05 6.30 ;
        RECT  12.55 2.45 13.05 5.40 ;
        RECT  13.20 4.90 13.70 7.25 ;
        RECT  12.85 4.90 13.75 6.30 ;
        RECT  14.15 6.75 14.95 10.55 ;
        RECT  15.05 3.80 15.55 5.40 ;
        RECT  12.55 4.90 15.55 5.40 ;
        RECT  15.55 2.45 16.25 4.50 ;
        RECT  15.05 3.80 16.25 4.50 ;
        RECT  16.85 6.75 17.65 10.55 ;
        RECT  11.45 6.75 17.80 7.25 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.68 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.95 ;
        PORT
        LAYER M1M ;
        RECT  0.25 2.80 1.15 3.70 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 10.40 1.15 11.00 ;
        RECT  1.80 7.90 2.65 11.00 ;
        RECT  5.95 9.95 6.65 11.00 ;
        RECT  7.45 7.15 8.20 11.00 ;
        RECT  10.10 7.10 10.90 11.00 ;
        RECT  12.80 7.70 13.60 11.00 ;
        RECT  15.50 7.75 16.30 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.60 2.00 2.30 2.85 ;
        RECT  4.85 2.00 5.70 4.45 ;
        RECT  7.70 2.00 8.40 3.25 ;
        RECT  11.00 2.00 11.70 4.50 ;
        RECT  14.20 2.00 14.45 4.45 ;
        RECT  13.70 2.80 14.45 4.45 ;
        RECT  14.20 2.00 14.90 3.30 ;
        RECT  13.70 2.80 14.90 3.30 ;
        RECT  17.05 2.00 17.75 4.50 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 4.40 0.95 9.50 ;
        RECT  0.45 6.95 1.15 9.50 ;
        RECT  1.60 3.75 2.15 4.95 ;
        RECT  0.45 4.40 2.15 4.95 ;
        RECT  1.60 3.75 2.35 4.50 ;
        RECT  0.45 4.40 2.35 4.50 ;
        RECT  3.15 2.50 3.90 4.55 ;
        RECT  3.00 5.85 3.50 7.45 ;
        RECT  0.45 6.95 3.50 7.45 ;
        RECT  3.00 5.85 3.70 6.55 ;
        RECT  3.35 2.50 3.90 5.40 ;
        RECT  3.35 4.90 4.65 5.40 ;
        RECT  4.15 4.90 4.65 8.70 ;
        RECT  3.30 8.00 4.65 8.70 ;
        RECT  5.10 7.70 5.15 10.35 ;
        RECT  4.45 9.15 5.15 10.35 ;
        RECT  5.10 7.70 5.60 9.65 ;
        RECT  4.45 9.15 5.60 9.65 ;
        RECT  5.15 6.55 5.90 7.25 ;
        RECT  4.15 6.75 5.90 7.25 ;
        RECT  6.35 2.55 7.05 3.25 ;
        RECT  6.50 2.55 7.00 8.20 ;
        RECT  5.10 7.70 7.00 8.20 ;
        RECT  6.50 2.55 7.05 4.95 ;
        RECT  6.50 4.45 9.00 4.95 ;
        RECT  8.30 4.45 9.00 5.20 ;
        RECT  9.05 5.85 9.55 10.55 ;
        RECT  8.75 7.05 9.55 10.55 ;
        RECT  9.50 3.55 10.30 4.30 ;
        RECT  9.80 3.55 10.30 6.35 ;
        RECT  9.80 5.65 11.20 6.35 ;
        RECT  9.05 5.85 11.20 6.35 ;
    END
END ITLCX12
MACRO ITLCX16
    CLASS CORE ;
    FOREIGN ITLCX16 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  14.35 6.80 15.15 10.55 ;
        RECT  15.75 2.45 16.45 4.60 ;
        RECT  15.95 2.45 16.45 5.40 ;
        RECT  17.05 6.80 17.85 10.55 ;
        RECT  18.45 2.45 19.20 5.40 ;
        RECT  19.90 6.80 20.70 10.55 ;
        RECT  21.15 2.45 21.90 5.40 ;
        RECT  21.25 2.45 21.90 6.30 ;
        RECT  21.25 5.40 22.15 6.30 ;
        RECT  21.65 2.45 21.90 7.30 ;
        RECT  15.95 4.90 21.90 5.40 ;
        RECT  21.65 5.40 22.15 7.30 ;
        RECT  14.35 6.80 23.40 7.30 ;
        RECT  22.60 6.80 23.40 10.55 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.73 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.50 2.55 7.60 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.33 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.20 8.30 3.00 11.00 ;
        RECT  3.70 7.20 4.50 11.00 ;
        RECT  7.65 7.40 8.40 11.00 ;
        RECT  10.30 7.70 11.10 11.00 ;
        RECT  13.00 7.75 13.80 11.00 ;
        RECT  15.70 7.75 16.50 11.00 ;
        RECT  18.45 7.75 19.30 11.00 ;
        RECT  21.25 7.75 22.05 11.00 ;
        RECT  0.00 11.00 23.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.75 2.00 2.55 2.90 ;
        RECT  5.35 2.00 6.05 4.40 ;
        RECT  5.35 2.00 7.25 2.25 ;
        RECT  9.25 2.00 9.95 4.00 ;
        RECT  11.00 2.00 13.55 2.10 ;
        RECT  14.40 2.00 15.10 4.50 ;
        RECT  17.10 2.00 17.80 4.45 ;
        RECT  19.80 2.00 20.50 4.45 ;
        RECT  22.65 2.00 23.35 4.50 ;
        RECT  0.00 0.00 23.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.70 5.55 1.20 10.55 ;
        RECT  0.70 8.30 1.65 10.55 ;
        RECT  1.85 3.55 2.35 6.05 ;
        RECT  1.75 3.55 2.45 4.25 ;
        RECT  0.70 5.55 3.70 6.05 ;
        RECT  3.50 2.50 4.20 3.20 ;
        RECT  3.00 5.40 3.70 6.10 ;
        RECT  3.70 2.50 4.20 4.25 ;
        RECT  3.70 3.55 4.90 4.25 ;
        RECT  4.40 3.55 4.90 5.35 ;
        RECT  4.40 4.85 5.45 5.35 ;
        RECT  4.95 4.85 5.45 10.55 ;
        RECT  4.95 9.85 7.10 10.55 ;
        RECT  6.70 2.80 7.20 8.85 ;
        RECT  6.05 7.25 7.20 8.85 ;
        RECT  6.70 2.80 7.40 4.95 ;
        RECT  7.90 2.55 8.60 3.30 ;
        RECT  6.70 2.80 8.60 3.30 ;
        RECT  8.95 6.75 9.75 10.55 ;
        RECT  6.70 4.45 12.85 4.95 ;
        RECT  11.75 3.30 12.45 4.00 ;
        RECT  12.00 5.85 12.45 10.55 ;
        RECT  11.65 6.75 12.45 10.55 ;
        RECT  12.00 5.85 12.50 7.25 ;
        RECT  8.95 6.75 12.50 7.25 ;
        RECT  12.15 4.45 12.85 5.15 ;
        RECT  11.75 3.50 13.95 4.00 ;
        RECT  13.45 3.50 13.95 6.35 ;
        RECT  13.45 5.65 14.20 6.35 ;
        RECT  12.00 5.85 14.20 6.35 ;
    END
END ITLCX16
MACRO ITLCX20
    CLASS CORE ;
    FOREIGN ITLCX20 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 25.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  14.35 6.80 15.15 10.55 ;
        RECT  15.75 2.45 16.45 4.60 ;
        RECT  15.95 2.45 16.45 5.40 ;
        RECT  17.05 6.80 17.85 10.55 ;
        RECT  18.45 2.45 19.20 5.40 ;
        RECT  19.75 6.80 20.55 10.55 ;
        RECT  21.15 2.45 21.90 5.40 ;
        RECT  21.25 2.45 21.90 6.30 ;
        RECT  21.25 5.40 22.15 6.30 ;
        RECT  21.65 2.45 21.90 7.30 ;
        RECT  15.95 4.90 21.90 5.40 ;
        RECT  21.65 5.40 22.15 7.30 ;
        RECT  14.35 6.80 23.25 7.30 ;
        RECT  22.45 6.80 23.25 10.55 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.73 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.50 2.55 7.60 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.33 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.20 8.30 3.00 11.00 ;
        RECT  3.75 7.20 4.45 11.00 ;
        RECT  7.65 7.40 8.40 11.00 ;
        RECT  10.30 7.70 11.10 11.00 ;
        RECT  13.00 7.75 13.80 11.00 ;
        RECT  15.70 7.75 16.50 11.00 ;
        RECT  18.45 7.75 19.15 11.00 ;
        RECT  21.10 7.75 21.90 11.00 ;
        RECT  23.95 6.90 24.75 11.00 ;
        RECT  0.00 11.00 25.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.60 2.00 2.40 2.90 ;
        RECT  5.35 2.00 6.05 4.40 ;
        RECT  5.35 2.00 7.25 2.25 ;
        RECT  9.25 2.00 9.95 4.00 ;
        RECT  11.00 2.00 13.55 2.10 ;
        RECT  14.40 2.00 15.10 4.50 ;
        RECT  17.10 2.00 17.80 4.45 ;
        RECT  19.80 2.00 20.50 4.45 ;
        RECT  22.50 2.00 23.20 4.55 ;
        RECT  24.05 2.00 24.75 4.50 ;
        RECT  0.00 0.00 25.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.70 5.55 1.20 10.55 ;
        RECT  0.70 8.25 1.65 10.55 ;
        RECT  1.60 3.55 2.10 6.05 ;
        RECT  1.60 3.55 2.30 4.25 ;
        RECT  0.70 5.55 3.75 6.05 ;
        RECT  3.50 2.45 4.20 3.15 ;
        RECT  3.05 5.40 3.75 6.10 ;
        RECT  3.70 2.45 4.20 4.25 ;
        RECT  3.70 3.55 4.90 4.25 ;
        RECT  4.40 3.55 4.90 5.45 ;
        RECT  4.40 4.85 5.45 5.45 ;
        RECT  4.95 4.85 5.45 10.55 ;
        RECT  4.95 9.80 7.15 10.55 ;
        RECT  6.70 2.80 7.20 8.85 ;
        RECT  6.05 7.25 7.20 8.85 ;
        RECT  6.70 2.80 7.40 4.95 ;
        RECT  7.90 2.55 8.60 3.30 ;
        RECT  6.70 2.80 8.60 3.30 ;
        RECT  8.95 6.75 9.75 10.55 ;
        RECT  6.70 4.45 12.85 4.95 ;
        RECT  11.75 3.30 12.45 4.00 ;
        RECT  12.00 5.85 12.45 10.55 ;
        RECT  11.65 6.75 12.45 10.55 ;
        RECT  12.00 5.85 12.50 7.25 ;
        RECT  8.95 6.75 12.50 7.25 ;
        RECT  12.15 4.45 12.85 5.15 ;
        RECT  11.75 3.50 13.95 4.00 ;
        RECT  13.45 3.50 13.95 6.35 ;
        RECT  13.45 5.65 14.20 6.35 ;
        RECT  12.00 5.85 14.20 6.35 ;
    END
END ITLCX20
MACRO ITLCX3
    CLASS CORE ;
    FOREIGN ITLCX3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.30 6.75 10.80 10.55 ;
        RECT  10.00 7.95 10.80 10.55 ;
        RECT  11.40 2.45 12.10 4.60 ;
        RECT  11.65 2.45 12.10 7.25 ;
        RECT  11.60 2.45 12.10 6.30 ;
        RECT  11.65 5.40 12.15 7.25 ;
        RECT  10.30 6.75 12.15 7.25 ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.16 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.55 7.60 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.67 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 8.05 2.70 11.00 ;
        RECT  1.85 10.10 4.05 11.00 ;
        RECT  0.40 10.85 4.05 11.00 ;
        RECT  5.95 9.20 6.75 11.00 ;
        RECT  4.85 9.70 6.75 11.00 ;
        RECT  8.65 9.05 9.45 11.00 ;
        RECT  11.35 7.95 12.15 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  4.15 2.00 4.95 4.25 ;
        RECT  6.85 2.00 7.65 4.40 ;
        RECT  10.05 2.00 10.75 4.50 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.25 5.65 0.75 9.75 ;
        RECT  0.25 8.75 1.20 9.75 ;
        RECT  0.90 2.95 2.10 3.65 ;
        RECT  1.60 2.95 2.10 6.15 ;
        RECT  2.55 2.45 3.25 4.50 ;
        RECT  0.25 5.65 3.65 6.15 ;
        RECT  2.75 2.45 3.25 5.20 ;
        RECT  2.95 5.65 3.65 6.35 ;
        RECT  2.75 4.70 4.60 5.20 ;
        RECT  4.10 4.70 4.60 8.75 ;
        RECT  3.35 7.75 4.60 8.75 ;
        RECT  5.45 3.50 5.95 7.80 ;
        RECT  5.05 7.10 5.95 7.80 ;
        RECT  5.45 3.50 6.25 5.55 ;
        RECT  6.40 6.90 6.90 8.75 ;
        RECT  3.35 8.25 6.90 8.75 ;
        RECT  6.40 6.90 7.60 7.60 ;
        RECT  7.30 4.85 8.00 5.55 ;
        RECT  5.45 5.05 8.00 5.55 ;
        RECT  7.60 8.10 8.10 10.55 ;
        RECT  7.35 8.95 8.10 10.55 ;
        RECT  8.50 3.70 9.30 4.45 ;
        RECT  8.80 3.70 9.30 8.60 ;
        RECT  7.60 8.10 9.30 8.60 ;
        RECT  8.80 6.80 9.85 7.50 ;
    END
END ITLCX3
MACRO ITLCX4
    CLASS CORE ;
    FOREIGN ITLCX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.30 6.75 10.80 10.55 ;
        RECT  10.00 7.95 10.80 10.55 ;
        RECT  11.25 2.45 11.95 4.60 ;
        RECT  11.65 2.45 11.95 7.25 ;
        RECT  11.45 2.45 11.95 6.30 ;
        RECT  11.65 5.40 12.15 7.25 ;
        RECT  10.30 6.75 12.15 7.25 ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.16 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.55 7.60 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.67 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 8.05 2.70 11.00 ;
        RECT  1.85 10.10 4.05 11.00 ;
        RECT  0.40 10.85 4.05 11.00 ;
        RECT  5.95 9.20 6.75 11.00 ;
        RECT  4.85 9.70 6.75 11.00 ;
        RECT  8.65 9.05 9.45 11.00 ;
        RECT  11.35 7.95 12.15 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  4.15 2.00 4.95 4.25 ;
        RECT  6.85 2.00 7.65 4.40 ;
        RECT  9.90 2.00 10.60 4.50 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.25 5.65 0.75 9.75 ;
        RECT  0.25 8.75 1.20 9.75 ;
        RECT  0.90 2.95 2.10 3.65 ;
        RECT  1.60 2.95 2.10 6.15 ;
        RECT  2.55 2.45 3.25 4.50 ;
        RECT  0.25 5.65 3.65 6.15 ;
        RECT  2.75 2.45 3.25 5.20 ;
        RECT  2.95 5.65 3.65 6.35 ;
        RECT  2.75 4.70 4.60 5.20 ;
        RECT  4.10 4.70 4.60 8.75 ;
        RECT  3.35 7.75 4.60 8.75 ;
        RECT  5.45 3.50 5.95 7.80 ;
        RECT  5.05 7.10 5.95 7.80 ;
        RECT  5.45 3.50 6.25 5.55 ;
        RECT  6.40 6.90 6.90 8.75 ;
        RECT  3.35 8.25 6.90 8.75 ;
        RECT  6.40 6.90 7.60 7.60 ;
        RECT  7.30 4.85 8.00 5.55 ;
        RECT  5.45 5.05 8.00 5.55 ;
        RECT  7.60 8.10 8.10 10.55 ;
        RECT  7.35 8.95 8.10 10.55 ;
        RECT  8.35 3.70 9.30 4.45 ;
        RECT  8.80 3.70 9.30 8.60 ;
        RECT  7.60 8.10 9.30 8.60 ;
        RECT  8.80 6.80 9.85 7.50 ;
    END
END ITLCX4
MACRO ITLCX8
    CLASS CORE ;
    FOREIGN ITLCX8 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.45 6.75 12.25 10.55 ;
        RECT  12.40 2.45 13.10 4.60 ;
        RECT  12.60 2.45 13.10 6.30 ;
        RECT  13.20 5.40 13.70 7.25 ;
        RECT  12.60 5.40 13.75 6.30 ;
        RECT  11.45 6.75 14.95 7.25 ;
        RECT  14.15 6.75 14.95 10.55 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.68 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.95 ;
        PORT
        LAYER M1M ;
        RECT  0.25 2.80 1.15 3.70 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 10.40 1.15 11.00 ;
        RECT  1.80 7.90 2.65 11.00 ;
        RECT  5.95 9.95 6.65 11.00 ;
        RECT  7.45 7.70 8.20 11.00 ;
        RECT  10.10 7.10 10.90 11.00 ;
        RECT  12.80 7.70 13.60 11.00 ;
        RECT  15.50 7.15 16.30 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.60 2.00 2.30 2.85 ;
        RECT  4.85 2.00 5.70 4.45 ;
        RECT  7.70 2.00 8.40 3.25 ;
        RECT  11.05 2.00 11.75 4.50 ;
        RECT  14.10 2.00 14.85 4.45 ;
        RECT  13.75 3.40 14.85 4.45 ;
        RECT  15.65 2.00 16.35 4.50 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 4.40 0.95 9.50 ;
        RECT  0.45 6.95 1.15 9.50 ;
        RECT  1.60 3.75 2.15 4.95 ;
        RECT  0.45 4.40 2.15 4.95 ;
        RECT  1.60 3.75 2.35 4.50 ;
        RECT  0.45 4.40 2.35 4.50 ;
        RECT  3.15 2.50 3.90 4.55 ;
        RECT  3.00 5.85 3.50 7.45 ;
        RECT  0.45 6.95 3.50 7.45 ;
        RECT  3.00 5.85 3.70 6.55 ;
        RECT  3.35 2.50 3.90 5.40 ;
        RECT  3.35 4.90 4.65 5.40 ;
        RECT  4.15 4.90 4.65 8.70 ;
        RECT  3.30 8.00 4.65 8.70 ;
        RECT  5.10 7.70 5.15 10.35 ;
        RECT  4.45 9.15 5.15 10.35 ;
        RECT  5.10 7.70 5.60 9.65 ;
        RECT  4.45 9.15 5.60 9.65 ;
        RECT  5.15 6.55 5.90 7.25 ;
        RECT  4.15 6.75 5.90 7.25 ;
        RECT  6.35 2.55 7.05 3.25 ;
        RECT  6.50 2.55 7.00 8.20 ;
        RECT  5.10 7.70 7.00 8.20 ;
        RECT  6.50 2.55 7.05 4.95 ;
        RECT  6.50 4.45 9.10 4.95 ;
        RECT  8.40 4.45 9.10 5.20 ;
        RECT  9.05 5.85 9.55 10.55 ;
        RECT  8.75 7.05 9.55 10.55 ;
        RECT  9.55 3.55 10.30 4.30 ;
        RECT  9.80 3.55 10.30 6.35 ;
        RECT  9.80 5.65 11.20 6.35 ;
        RECT  9.05 5.85 11.20 6.35 ;
    END
END ITLCX8
MACRO ITLX1
    CLASS CORE ;
    FOREIGN ITLX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.30 2.70 5.35 4.40 ;
        RECT  4.85 2.70 5.35 10.55 ;
        RECT  4.30 7.70 5.35 10.55 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  0.25 9.30 1.15 10.20 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 3.10 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.95 7.70 2.65 11.00 ;
        RECT  0.00 11.00 5.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.95 2.00 2.65 4.45 ;
        RECT  0.00 0.00 5.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.75 0.95 8.85 ;
        RECT  0.45 3.75 1.15 4.45 ;
        RECT  0.45 6.75 1.15 8.85 ;
        RECT  3.65 4.85 4.15 7.25 ;
        RECT  0.45 6.75 4.15 7.25 ;
        RECT  3.65 4.85 4.35 5.55 ;
    END
END ITLX1
MACRO ITLX12
    CLASS CORE ;
    FOREIGN ITLX12 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.65 8.00 9.55 8.90 ;
        RECT  8.80 2.45 9.55 4.05 ;
        RECT  9.00 2.45 9.55 10.55 ;
        RECT  8.80 7.70 9.55 10.55 ;
        RECT  11.50 6.50 12.00 10.55 ;
        RECT  11.50 2.45 12.20 4.90 ;
        RECT  11.50 7.70 12.20 10.55 ;
        RECT  9.00 6.50 14.70 7.00 ;
        RECT  14.20 2.45 14.70 4.90 ;
        RECT  9.00 4.40 14.70 4.90 ;
        RECT  14.20 6.50 14.70 10.55 ;
        RECT  14.20 2.45 14.90 4.05 ;
        RECT  14.20 7.70 14.90 10.55 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.65 9.25 1.35 11.00 ;
        RECT  4.60 9.95 5.30 11.00 ;
        RECT  7.45 7.70 8.15 11.00 ;
        RECT  10.15 7.55 10.85 11.00 ;
        RECT  12.85 7.55 13.55 11.00 ;
        RECT  15.55 7.70 16.25 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.60 ;
        RECT  7.45 2.00 8.15 4.00 ;
        RECT  10.15 2.00 10.85 3.95 ;
        RECT  12.85 2.00 13.55 3.95 ;
        RECT  15.55 2.00 16.25 4.00 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.80 6.85 3.95 7.35 ;
        RECT  1.60 7.75 2.50 8.25 ;
        RECT  0.95 3.25 2.10 3.95 ;
        RECT  1.40 3.25 2.10 5.00 ;
        RECT  2.00 3.25 2.10 10.55 ;
        RECT  1.60 3.25 2.10 8.25 ;
        RECT  2.00 7.75 2.50 10.55 ;
        RECT  2.55 3.45 3.30 4.15 ;
        RECT  3.25 3.45 3.30 9.40 ;
        RECT  2.80 3.45 3.30 7.35 ;
        RECT  3.25 6.85 3.95 9.40 ;
        RECT  2.00 9.85 4.15 10.55 ;
        RECT  4.10 2.55 4.80 4.95 ;
        RECT  4.80 4.45 5.30 8.45 ;
        RECT  4.60 6.85 5.30 8.45 ;
        RECT  3.25 8.90 6.80 9.40 ;
        RECT  6.10 2.45 6.80 4.95 ;
        RECT  6.30 6.75 6.80 10.55 ;
        RECT  6.10 7.70 6.80 10.55 ;
        RECT  4.10 4.45 8.50 4.95 ;
        RECT  7.80 4.45 8.50 5.15 ;
        RECT  7.85 6.50 8.55 7.25 ;
        RECT  6.30 6.75 8.55 7.25 ;
        RECT  10.00 5.35 10.70 6.05 ;
        RECT  10.00 5.55 16.60 6.05 ;
        RECT  16.10 4.45 16.60 7.25 ;
        RECT  16.10 6.75 17.55 7.25 ;
        RECT  17.05 3.35 17.55 4.95 ;
        RECT  16.10 4.45 17.55 4.95 ;
        RECT  17.05 6.75 17.55 9.40 ;
        RECT  17.05 3.35 17.75 4.05 ;
        RECT  17.05 7.70 17.75 9.40 ;
    END
END ITLX12
MACRO ITLX16
    CLASS CORE ;
    FOREIGN ITLX16 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.65 2.80 9.60 3.70 ;
        RECT  8.90 2.45 9.60 4.05 ;
        RECT  9.30 2.45 9.60 10.55 ;
        RECT  9.10 2.45 9.60 4.90 ;
        RECT  9.30 4.40 9.80 10.55 ;
        RECT  9.00 7.70 9.80 10.55 ;
        RECT  11.60 2.45 12.30 4.90 ;
        RECT  11.70 6.50 12.40 10.55 ;
        RECT  14.30 2.45 15.00 4.90 ;
        RECT  14.40 6.50 15.10 10.55 ;
        RECT  9.30 6.50 17.60 7.00 ;
        RECT  17.00 2.45 17.50 4.90 ;
        RECT  9.10 4.40 17.50 4.90 ;
        RECT  17.10 6.50 17.60 10.55 ;
        RECT  17.00 2.45 17.70 4.05 ;
        RECT  17.10 7.70 17.80 10.55 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.65 9.25 1.35 11.00 ;
        RECT  4.35 9.95 5.05 11.00 ;
        RECT  7.65 7.70 8.35 11.00 ;
        RECT  10.35 7.55 11.05 11.00 ;
        RECT  13.05 7.55 13.75 11.00 ;
        RECT  15.75 7.55 16.45 11.00 ;
        RECT  18.45 7.70 19.15 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.60 ;
        RECT  7.40 2.00 8.10 4.00 ;
        RECT  10.25 2.00 10.95 3.95 ;
        RECT  12.95 2.00 13.65 3.95 ;
        RECT  15.65 2.00 16.35 3.95 ;
        RECT  18.35 2.00 19.05 4.00 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.80 6.85 3.70 7.35 ;
        RECT  1.60 7.85 2.50 8.35 ;
        RECT  0.95 3.25 2.10 3.95 ;
        RECT  1.40 3.25 2.10 5.00 ;
        RECT  2.00 3.25 2.10 10.55 ;
        RECT  1.60 3.25 2.10 8.35 ;
        RECT  2.00 7.85 2.50 10.55 ;
        RECT  2.55 3.45 3.30 4.15 ;
        RECT  3.00 3.45 3.30 9.40 ;
        RECT  2.80 3.45 3.30 7.35 ;
        RECT  3.00 6.85 3.70 9.40 ;
        RECT  2.00 9.85 3.90 10.55 ;
        RECT  4.55 2.55 4.80 8.45 ;
        RECT  4.10 2.55 4.80 4.95 ;
        RECT  4.55 4.45 5.05 8.45 ;
        RECT  4.35 6.85 5.05 8.45 ;
        RECT  3.00 8.90 6.75 9.40 ;
        RECT  6.05 2.45 6.75 4.95 ;
        RECT  6.40 6.75 6.75 10.55 ;
        RECT  6.05 8.05 6.75 10.55 ;
        RECT  6.40 6.75 6.90 9.00 ;
        RECT  3.00 8.90 6.90 9.00 ;
        RECT  4.10 4.45 8.65 4.95 ;
        RECT  7.95 4.45 8.65 5.15 ;
        RECT  8.15 6.50 8.85 7.25 ;
        RECT  6.40 6.75 8.85 7.25 ;
        RECT  10.25 5.35 10.95 6.05 ;
        RECT  10.25 5.55 19.40 6.05 ;
        RECT  18.90 4.45 19.40 7.25 ;
        RECT  18.90 6.75 20.35 7.25 ;
        RECT  19.85 3.35 20.35 4.95 ;
        RECT  18.90 4.45 20.35 4.95 ;
        RECT  19.85 6.75 20.35 9.40 ;
        RECT  19.85 3.35 20.55 4.05 ;
        RECT  19.85 7.70 20.55 9.40 ;
    END
END ITLX16
MACRO ITLX2
    CLASS CORE ;
    FOREIGN ITLX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.80 2.45 9.30 10.55 ;
        RECT  8.60 7.80 9.30 10.55 ;
        RECT  8.65 2.45 9.55 4.05 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.45 1.15 11.00 ;
        RECT  4.40 10.25 5.10 11.00 ;
        RECT  7.25 7.80 7.95 11.00 ;
        RECT  11.45 7.15 12.15 11.00 ;
        RECT  10.25 10.10 12.15 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.75 ;
        RECT  7.35 2.00 8.05 4.00 ;
        RECT  10.40 2.00 11.10 3.15 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.65 4.70 2.35 5.40 ;
        RECT  2.80 5.40 3.80 5.90 ;
        RECT  0.95 3.40 2.15 4.10 ;
        RECT  1.80 3.40 2.15 10.25 ;
        RECT  1.65 3.40 2.15 5.40 ;
        RECT  1.80 4.70 2.35 10.25 ;
        RECT  1.80 7.45 2.50 10.25 ;
        RECT  2.60 3.60 3.30 4.30 ;
        RECT  1.80 9.55 2.85 10.25 ;
        RECT  2.80 3.60 3.30 5.90 ;
        RECT  3.30 5.40 3.80 9.80 ;
        RECT  3.30 7.15 4.00 9.80 ;
        RECT  4.65 2.70 4.85 8.85 ;
        RECT  4.15 2.70 4.85 4.95 ;
        RECT  4.65 4.45 5.15 8.85 ;
        RECT  4.65 7.15 5.35 8.85 ;
        RECT  3.30 9.30 6.45 9.80 ;
        RECT  5.95 6.85 6.45 10.55 ;
        RECT  5.75 9.30 6.45 10.55 ;
        RECT  5.85 3.35 6.55 4.95 ;
        RECT  4.15 4.45 8.35 4.95 ;
        RECT  7.65 4.45 8.35 5.15 ;
        RECT  7.65 6.65 8.35 7.35 ;
        RECT  5.95 6.85 8.35 7.35 ;
        RECT  9.75 5.85 10.80 6.55 ;
        RECT  10.30 3.80 10.80 8.85 ;
        RECT  10.10 5.85 10.80 8.85 ;
        RECT  10.30 3.80 11.10 4.50 ;
    END
END ITLX2
MACRO ITLX20
    CLASS CORE ;
    FOREIGN ITLX20 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  9.00 2.45 9.75 4.05 ;
        RECT  9.55 2.45 9.75 10.55 ;
        RECT  9.25 2.45 9.75 4.90 ;
        RECT  9.55 4.40 10.05 10.55 ;
        RECT  9.15 7.75 10.05 10.55 ;
        RECT  11.70 2.45 12.40 4.90 ;
        RECT  11.85 6.50 12.55 10.55 ;
        RECT  14.40 2.45 15.10 4.90 ;
        RECT  14.55 6.50 15.25 10.55 ;
        RECT  17.05 6.50 17.95 7.60 ;
        RECT  17.10 2.45 17.80 4.90 ;
        RECT  17.25 6.50 17.95 10.55 ;
        RECT  9.55 6.50 20.65 7.00 ;
        RECT  19.80 2.45 20.50 4.90 ;
        RECT  9.25 4.40 20.50 4.90 ;
        RECT  19.95 6.50 20.65 10.55 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  22.65 5.40 23.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 9.90 1.15 11.00 ;
        RECT  3.35 9.95 4.05 11.00 ;
        RECT  7.75 7.75 8.45 11.00 ;
        RECT  10.50 7.45 11.20 11.00 ;
        RECT  13.20 7.45 13.90 11.00 ;
        RECT  15.90 7.45 16.60 11.00 ;
        RECT  18.60 7.45 19.30 11.00 ;
        RECT  21.30 7.70 22.00 11.00 ;
        RECT  0.00 11.00 23.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.50 ;
        RECT  7.65 2.00 8.35 4.00 ;
        RECT  10.35 2.00 11.05 3.95 ;
        RECT  13.05 2.00 13.75 3.95 ;
        RECT  15.75 2.00 16.45 3.95 ;
        RECT  18.45 2.00 19.15 3.95 ;
        RECT  21.15 2.00 21.85 4.00 ;
        RECT  0.00 0.00 23.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.95 4.20 2.10 4.90 ;
        RECT  1.40 8.00 2.10 8.70 ;
        RECT  1.60 3.15 1.65 10.55 ;
        RECT  0.95 3.15 1.65 4.90 ;
        RECT  1.60 4.20 2.10 10.55 ;
        RECT  1.60 9.85 2.50 10.55 ;
        RECT  2.50 3.05 3.30 3.75 ;
        RECT  2.55 6.45 3.30 8.05 ;
        RECT  2.80 3.05 3.30 9.50 ;
        RECT  4.05 2.45 4.60 8.20 ;
        RECT  3.90 6.50 4.60 8.20 ;
        RECT  2.80 9.00 5.20 9.50 ;
        RECT  4.05 2.45 4.75 4.95 ;
        RECT  4.70 9.00 5.20 10.55 ;
        RECT  5.85 2.45 7.00 3.15 ;
        RECT  5.45 7.90 7.00 8.60 ;
        RECT  6.30 7.90 7.00 10.55 ;
        RECT  6.30 2.45 7.00 4.95 ;
        RECT  6.50 6.80 7.00 10.55 ;
        RECT  4.70 9.85 7.00 10.55 ;
        RECT  4.05 4.45 8.75 4.95 ;
        RECT  8.05 4.45 8.75 5.25 ;
        RECT  8.35 6.60 9.10 7.30 ;
        RECT  6.50 6.80 9.10 7.30 ;
        RECT  10.50 5.35 11.20 6.05 ;
        RECT  10.50 5.55 22.20 6.05 ;
        RECT  21.70 4.45 22.20 7.25 ;
        RECT  21.70 6.75 23.15 7.25 ;
        RECT  22.65 3.35 23.15 4.95 ;
        RECT  21.70 4.45 23.15 4.95 ;
        RECT  22.65 6.75 23.15 9.40 ;
        RECT  22.65 3.35 23.35 4.05 ;
        RECT  22.65 7.70 23.35 9.40 ;
    END
END ITLX20
MACRO ITLX3
    CLASS CORE ;
    FOREIGN ITLX3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.80 2.80 9.30 10.20 ;
        RECT  8.60 7.60 9.35 10.20 ;
        RECT  8.65 2.80 9.55 3.70 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  10.05 4.10 11.20 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.15 1.15 11.00 ;
        RECT  4.40 10.25 5.10 11.00 ;
        RECT  7.25 7.70 7.95 11.00 ;
        RECT  7.10 9.75 7.95 11.00 ;
        RECT  9.95 7.40 10.65 11.00 ;
        RECT  9.95 10.10 12.15 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 3.00 ;
        RECT  7.35 2.00 8.05 3.55 ;
        RECT  10.05 2.00 10.75 3.30 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.65 4.70 2.35 5.40 ;
        RECT  2.80 5.40 3.80 5.90 ;
        RECT  1.80 3.65 2.15 8.85 ;
        RECT  1.80 7.15 2.50 8.85 ;
        RECT  0.95 3.65 2.15 4.35 ;
        RECT  2.00 3.65 2.15 10.55 ;
        RECT  1.65 3.65 2.15 5.40 ;
        RECT  2.00 4.70 2.35 10.55 ;
        RECT  1.80 4.70 2.35 8.85 ;
        RECT  2.00 7.15 2.50 10.55 ;
        RECT  2.60 3.60 3.30 4.30 ;
        RECT  2.00 9.85 2.85 10.55 ;
        RECT  2.80 3.60 3.30 5.90 ;
        RECT  3.30 5.40 3.80 9.80 ;
        RECT  3.30 7.15 4.00 9.80 ;
        RECT  4.65 2.70 4.85 8.85 ;
        RECT  4.15 2.70 4.85 4.70 ;
        RECT  4.65 4.20 5.15 8.85 ;
        RECT  4.65 7.15 5.35 8.85 ;
        RECT  3.30 9.30 6.45 9.80 ;
        RECT  5.95 6.45 6.45 10.55 ;
        RECT  5.75 9.30 6.45 10.55 ;
        RECT  5.85 3.10 6.55 4.70 ;
        RECT  4.15 4.20 8.35 4.70 ;
        RECT  7.65 4.20 8.35 4.90 ;
        RECT  7.65 6.25 8.35 6.95 ;
        RECT  5.95 6.45 8.35 6.95 ;
        RECT  9.75 5.45 10.45 6.15 ;
        RECT  11.45 2.60 12.15 3.30 ;
        RECT  9.75 5.45 12.15 5.95 ;
        RECT  11.65 2.60 12.15 9.00 ;
        RECT  11.45 7.40 12.15 9.00 ;
    END
END ITLX3
MACRO ITLX4
    CLASS CORE ;
    FOREIGN ITLX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.60 2.45 9.30 4.05 ;
        RECT  8.80 2.45 9.30 10.55 ;
        RECT  8.60 7.70 9.30 10.55 ;
        RECT  8.60 7.70 9.55 8.90 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  11.45 9.30 12.35 10.20 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.45 1.15 11.00 ;
        RECT  4.40 10.25 5.10 11.00 ;
        RECT  7.25 7.70 7.95 11.00 ;
        RECT  10.10 7.25 10.80 11.00 ;
        RECT  9.95 9.75 10.80 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.75 ;
        RECT  7.25 2.00 7.95 4.00 ;
        RECT  9.95 2.00 10.65 4.00 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.45 4.55 2.65 5.05 ;
        RECT  3.10 7.15 4.00 8.90 ;
        RECT  0.95 3.40 1.95 4.10 ;
        RECT  1.80 3.40 1.95 10.55 ;
        RECT  1.45 3.40 1.95 5.05 ;
        RECT  1.80 4.55 2.30 10.55 ;
        RECT  1.80 7.40 2.50 10.55 ;
        RECT  1.80 4.55 2.65 5.25 ;
        RECT  1.80 9.85 2.85 10.55 ;
        RECT  2.50 3.40 3.60 4.10 ;
        RECT  3.50 3.40 3.60 9.80 ;
        RECT  3.10 3.40 3.60 8.90 ;
        RECT  3.50 7.15 4.00 9.80 ;
        RECT  4.65 2.55 4.75 8.85 ;
        RECT  4.05 2.55 4.75 4.95 ;
        RECT  4.65 4.45 5.20 8.85 ;
        RECT  4.65 7.15 5.35 8.85 ;
        RECT  3.50 9.30 6.45 9.80 ;
        RECT  5.75 3.35 6.45 4.95 ;
        RECT  5.95 6.75 6.45 10.55 ;
        RECT  5.75 9.30 6.45 10.55 ;
        RECT  4.05 4.45 8.35 4.95 ;
        RECT  7.65 4.45 8.35 5.15 ;
        RECT  7.65 6.55 8.35 7.25 ;
        RECT  5.95 6.75 8.35 7.25 ;
        RECT  9.75 5.25 11.95 5.95 ;
        RECT  11.45 3.35 11.95 8.85 ;
        RECT  11.45 3.35 12.15 4.05 ;
        RECT  11.45 7.25 12.15 8.85 ;
    END
END ITLX4
MACRO ITLX8
    CLASS CORE ;
    FOREIGN ITLX8 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.65 2.45 9.55 4.05 ;
        RECT  9.05 2.45 9.55 10.55 ;
        RECT  8.80 7.70 9.55 10.55 ;
        RECT  9.05 6.55 11.90 7.05 ;
        RECT  11.40 2.45 11.90 4.90 ;
        RECT  9.05 4.40 11.90 4.90 ;
        RECT  11.40 6.55 11.90 10.55 ;
        RECT  11.40 2.45 12.10 4.05 ;
        RECT  11.40 7.70 12.20 10.55 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.65 9.25 1.35 11.00 ;
        RECT  4.60 9.95 5.30 11.00 ;
        RECT  7.45 7.70 8.15 11.00 ;
        RECT  10.15 7.55 10.85 11.00 ;
        RECT  12.85 7.70 13.55 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.60 ;
        RECT  7.35 2.00 8.05 4.00 ;
        RECT  10.05 2.00 10.75 3.95 ;
        RECT  12.75 2.00 13.45 4.00 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.80 6.85 3.95 7.35 ;
        RECT  1.60 7.80 2.50 8.30 ;
        RECT  0.95 3.25 2.10 3.95 ;
        RECT  1.40 3.25 2.10 5.00 ;
        RECT  2.00 3.25 2.10 10.55 ;
        RECT  1.60 3.25 2.10 8.30 ;
        RECT  2.00 7.80 2.50 10.55 ;
        RECT  2.55 3.45 3.30 4.15 ;
        RECT  3.25 3.45 3.30 9.40 ;
        RECT  2.80 3.45 3.30 7.35 ;
        RECT  3.25 6.85 3.95 9.40 ;
        RECT  2.00 9.85 4.15 10.55 ;
        RECT  4.10 2.55 4.80 4.95 ;
        RECT  4.80 4.45 5.30 8.45 ;
        RECT  4.60 6.85 5.30 8.45 ;
        RECT  3.25 8.90 6.80 9.40 ;
        RECT  6.00 2.45 6.70 4.95 ;
        RECT  6.30 6.75 6.80 10.55 ;
        RECT  6.10 7.70 6.80 10.55 ;
        RECT  4.10 4.45 8.40 4.95 ;
        RECT  7.70 4.45 8.40 5.15 ;
        RECT  7.90 6.50 8.60 7.25 ;
        RECT  6.30 6.75 8.60 7.25 ;
        RECT  10.00 5.35 10.70 6.05 ;
        RECT  10.00 5.55 13.80 6.05 ;
        RECT  13.30 4.45 13.80 7.25 ;
        RECT  13.30 6.75 14.75 7.25 ;
        RECT  14.25 3.35 14.75 4.95 ;
        RECT  13.30 4.45 14.75 4.95 ;
        RECT  14.25 6.75 14.75 9.40 ;
        RECT  14.25 3.35 14.95 4.05 ;
        RECT  14.25 7.70 14.95 9.40 ;
    END
END ITLX8
MACRO JKRRX1
    CLASS CORE ;
    FOREIGN JKRRX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 35.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  9.50 2.55 10.20 3.25 ;
        RECT  15.65 2.75 16.55 3.70 ;
        RECT  9.50 2.75 17.85 3.25 ;
        RECT  17.15 2.75 17.85 3.65 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M2M ;
        RECT  21.40 4.10 22.00 9.00 ;
        RECT  21.30 4.10 22.10 4.90 ;
        RECT  21.30 7.90 22.10 9.00 ;
        LAYER M1M ;
        RECT  21.35 8.00 22.05 9.75 ;
        RECT  21.25 8.00 22.15 8.90 ;
        RECT  21.55 3.75 22.25 4.95 ;
        RECT  21.25 4.05 22.25 4.95 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  24.25 3.75 24.95 4.45 ;
        RECT  24.45 3.75 24.75 9.75 ;
        RECT  24.05 7.95 24.75 9.75 ;
        RECT  24.45 3.75 24.95 8.95 ;
        RECT  24.05 7.95 24.95 8.95 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  26.85 4.10 27.75 5.00 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  33.85 5.40 34.75 6.30 ;
        END
    END J
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.25 6.65 2.55 7.35 ;
        RECT  1.65 6.65 2.55 7.65 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.30 2.50 11.00 ;
        RECT  4.05 7.95 4.75 11.00 ;
        RECT  9.80 8.20 10.50 11.00 ;
        RECT  12.30 9.55 13.00 11.00 ;
        RECT  17.15 9.05 17.85 11.00 ;
        RECT  19.85 9.15 20.55 11.00 ;
        RECT  22.70 8.25 23.40 11.00 ;
        RECT  27.55 8.50 28.25 11.00 ;
        RECT  32.40 10.65 33.10 11.00 ;
        RECT  0.00 11.00 35.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.90 2.00 1.70 3.20 ;
        RECT  4.05 2.00 4.75 4.85 ;
        RECT  2.70 2.00 5.20 2.50 ;
        RECT  8.50 2.00 9.00 4.25 ;
        RECT  9.90 3.75 10.60 4.95 ;
        RECT  8.50 3.75 13.60 4.25 ;
        RECT  12.90 3.75 13.60 5.40 ;
        RECT  18.30 2.00 18.35 5.40 ;
        RECT  17.60 4.65 18.35 5.40 ;
        RECT  18.30 2.00 18.80 5.15 ;
        RECT  17.60 4.65 18.80 5.15 ;
        RECT  18.30 2.00 21.75 2.90 ;
        RECT  22.90 2.00 23.60 4.40 ;
        RECT  22.90 2.00 25.55 2.55 ;
        RECT  26.55 2.00 27.25 3.65 ;
        RECT  31.25 2.00 31.95 3.65 ;
        RECT  0.00 0.00 35.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.25 5.35 0.75 10.25 ;
        RECT  0.25 9.55 1.15 10.25 ;
        RECT  1.00 3.80 1.80 5.85 ;
        RECT  0.25 5.35 1.80 5.85 ;
        RECT  2.70 4.20 3.55 4.90 ;
        RECT  3.05 4.20 3.55 8.85 ;
        RECT  2.70 8.15 3.55 8.85 ;
        RECT  3.05 5.55 6.35 6.05 ;
        RECT  5.35 3.20 5.85 6.05 ;
        RECT  5.85 5.55 6.35 7.40 ;
        RECT  5.85 6.70 6.55 7.40 ;
        RECT  6.40 4.20 7.55 4.90 ;
        RECT  6.85 3.00 7.55 3.70 ;
        RECT  5.35 3.20 7.55 3.70 ;
        RECT  7.05 4.20 7.55 9.25 ;
        RECT  6.40 8.55 8.00 9.25 ;
        RECT  9.35 5.65 10.05 6.35 ;
        RECT  10.35 6.90 11.05 7.60 ;
        RECT  7.05 7.10 11.05 7.60 ;
        RECT  11.40 4.75 12.10 6.15 ;
        RECT  9.35 5.65 12.10 6.15 ;
        RECT  11.60 4.75 12.10 8.85 ;
        RECT  11.15 8.10 12.10 8.85 ;
        RECT  15.25 4.70 15.50 9.85 ;
        RECT  14.80 7.15 15.50 9.85 ;
        RECT  15.25 4.70 15.75 7.65 ;
        RECT  15.25 4.70 15.95 5.40 ;
        RECT  16.95 5.95 17.65 6.70 ;
        RECT  18.50 8.15 19.20 9.85 ;
        RECT  19.00 6.95 19.70 7.65 ;
        RECT  14.80 7.15 19.70 7.65 ;
        RECT  20.00 4.75 20.70 6.45 ;
        RECT  16.95 5.95 20.70 6.45 ;
        RECT  20.20 4.75 20.70 8.65 ;
        RECT  18.50 8.15 20.70 8.65 ;
        RECT  20.00 5.75 23.95 6.25 ;
        RECT  23.25 5.55 23.95 6.25 ;
        RECT  16.95 5.95 23.95 6.25 ;
        RECT  25.45 6.45 26.15 7.20 ;
        RECT  25.50 5.25 26.20 5.95 ;
        RECT  26.55 7.50 27.05 9.25 ;
        RECT  26.20 7.65 27.05 9.25 ;
        RECT  26.55 7.50 29.60 8.00 ;
        RECT  26.20 7.65 29.60 8.00 ;
        RECT  28.90 2.95 29.60 4.80 ;
        RECT  28.90 7.50 29.60 9.15 ;
        RECT  29.80 9.65 30.50 10.35 ;
        RECT  30.25 6.45 30.95 8.15 ;
        RECT  30.60 5.25 31.30 5.95 ;
        RECT  25.50 5.45 31.30 5.95 ;
        RECT  28.90 4.30 32.30 4.80 ;
        RECT  31.60 7.50 32.10 9.15 ;
        RECT  28.90 8.65 32.10 9.15 ;
        RECT  31.80 4.30 32.30 6.95 ;
        RECT  25.45 6.45 32.30 6.95 ;
        RECT  31.60 7.50 32.30 8.25 ;
        RECT  32.60 2.95 33.30 3.65 ;
        RECT  32.80 2.95 33.30 10.15 ;
        RECT  29.80 9.65 34.45 10.15 ;
        RECT  33.75 9.65 34.45 10.35 ;
        LAYER V1M ;
        RECT  21.20 7.95 22.20 8.95 ;
        RECT  21.20 4.05 22.20 5.05 ;
    END
END JKRRX1
MACRO JKRRX2
    CLASS CORE ;
    FOREIGN JKRRX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 35.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  9.50 2.55 10.20 3.25 ;
        RECT  15.65 2.75 16.55 3.70 ;
        RECT  17.15 2.55 17.85 3.25 ;
        RECT  9.50 2.75 17.85 3.25 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M2M ;
        RECT  21.40 4.10 22.00 9.00 ;
        RECT  21.30 4.10 22.10 4.90 ;
        RECT  21.30 7.90 22.10 9.00 ;
        LAYER M1M ;
        RECT  21.35 7.85 22.05 10.55 ;
        RECT  21.25 7.85 22.15 8.90 ;
        RECT  21.55 2.75 22.25 4.95 ;
        RECT  21.25 4.05 22.25 4.95 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  24.25 2.75 24.95 4.45 ;
        RECT  24.45 2.75 24.75 10.55 ;
        RECT  24.05 7.85 24.75 10.55 ;
        RECT  24.45 2.75 24.95 8.95 ;
        RECT  24.05 7.85 24.95 8.95 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  26.85 4.10 27.75 5.00 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  33.85 5.40 34.75 6.30 ;
        END
    END J
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.25 6.65 2.55 7.35 ;
        RECT  1.65 6.65 2.55 7.65 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.30 2.50 11.00 ;
        RECT  4.05 7.95 4.75 11.00 ;
        RECT  9.80 8.20 10.50 11.00 ;
        RECT  12.30 9.55 13.00 11.00 ;
        RECT  17.15 9.05 17.85 11.00 ;
        RECT  19.85 9.15 20.55 11.00 ;
        RECT  22.70 7.90 23.40 11.00 ;
        RECT  27.55 8.50 28.25 11.00 ;
        RECT  32.40 10.65 33.10 11.00 ;
        RECT  0.00 11.00 35.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.90 2.00 1.70 3.20 ;
        RECT  4.05 2.00 4.75 4.85 ;
        RECT  2.70 2.00 5.20 2.50 ;
        RECT  8.50 2.00 9.00 4.25 ;
        RECT  9.90 3.75 10.60 4.95 ;
        RECT  8.50 3.75 13.60 4.25 ;
        RECT  12.90 3.75 13.60 5.00 ;
        RECT  18.30 2.00 18.35 5.00 ;
        RECT  17.60 4.25 18.35 5.00 ;
        RECT  18.30 2.00 18.80 4.75 ;
        RECT  17.60 4.25 18.80 4.75 ;
        RECT  22.90 2.00 23.60 4.40 ;
        RECT  26.55 2.00 27.25 3.65 ;
        RECT  31.25 2.00 31.95 3.65 ;
        RECT  0.00 0.00 35.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.25 5.35 0.75 10.25 ;
        RECT  0.25 9.55 1.15 10.25 ;
        RECT  1.00 3.80 1.80 5.85 ;
        RECT  0.25 5.35 1.80 5.85 ;
        RECT  2.70 4.20 3.55 4.90 ;
        RECT  3.05 4.20 3.55 8.85 ;
        RECT  2.70 8.15 3.55 8.85 ;
        RECT  3.05 5.55 6.35 6.05 ;
        RECT  5.35 3.20 5.85 6.05 ;
        RECT  5.85 5.55 6.35 7.40 ;
        RECT  5.85 6.70 6.55 7.40 ;
        RECT  6.40 4.20 7.55 4.90 ;
        RECT  6.85 3.00 7.55 3.70 ;
        RECT  5.35 3.20 7.55 3.70 ;
        RECT  7.05 4.20 7.55 9.25 ;
        RECT  6.40 8.55 8.00 9.25 ;
        RECT  9.35 5.65 10.05 6.35 ;
        RECT  10.35 6.90 11.05 7.60 ;
        RECT  7.05 7.10 11.05 7.60 ;
        RECT  11.40 4.75 12.10 6.15 ;
        RECT  9.35 5.65 12.10 6.15 ;
        RECT  11.60 4.75 12.10 8.85 ;
        RECT  11.15 8.10 12.10 8.85 ;
        RECT  15.25 4.30 15.50 9.85 ;
        RECT  14.80 7.15 15.50 9.85 ;
        RECT  15.25 4.30 15.75 7.65 ;
        RECT  15.25 4.30 15.95 5.00 ;
        RECT  16.95 5.95 17.65 6.70 ;
        RECT  18.50 8.15 19.20 9.85 ;
        RECT  19.00 6.95 19.70 7.65 ;
        RECT  14.80 7.15 19.70 7.65 ;
        RECT  20.00 4.35 20.70 6.45 ;
        RECT  16.95 5.95 20.70 6.45 ;
        RECT  20.20 4.35 20.70 8.65 ;
        RECT  18.50 8.15 20.70 8.65 ;
        RECT  20.00 5.75 23.95 6.25 ;
        RECT  23.25 5.55 23.95 6.25 ;
        RECT  16.95 5.95 23.95 6.25 ;
        RECT  25.45 6.45 26.15 7.20 ;
        RECT  25.50 5.25 26.20 5.95 ;
        RECT  26.55 7.50 27.05 9.25 ;
        RECT  26.20 7.65 27.05 9.25 ;
        RECT  26.55 7.50 29.60 8.00 ;
        RECT  26.20 7.65 29.60 8.00 ;
        RECT  28.90 2.95 29.60 4.80 ;
        RECT  28.90 7.50 29.60 9.15 ;
        RECT  29.80 9.65 30.50 10.35 ;
        RECT  30.25 6.45 30.95 8.15 ;
        RECT  30.60 5.25 31.30 5.95 ;
        RECT  25.50 5.45 31.30 5.95 ;
        RECT  28.90 4.30 32.30 4.80 ;
        RECT  31.60 7.50 32.10 9.15 ;
        RECT  28.90 8.65 32.10 9.15 ;
        RECT  31.80 4.30 32.30 6.95 ;
        RECT  25.45 6.45 32.30 6.95 ;
        RECT  31.60 7.50 32.30 8.25 ;
        RECT  32.60 2.95 33.30 3.65 ;
        RECT  32.80 2.95 33.30 10.15 ;
        RECT  29.80 9.65 34.45 10.15 ;
        RECT  33.75 9.65 34.45 10.35 ;
        LAYER V1M ;
        RECT  21.20 7.95 22.20 8.95 ;
        RECT  21.20 4.05 22.20 5.05 ;
    END
END JKRRX2
MACRO JKRRX4
    CLASS CORE ;
    FOREIGN JKRRX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 37.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  9.50 2.55 10.20 3.25 ;
        RECT  15.65 2.75 16.55 3.70 ;
        RECT  17.15 2.55 17.85 3.25 ;
        RECT  9.50 2.75 17.85 3.25 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M2M ;
        RECT  22.80 4.10 23.40 9.00 ;
        RECT  22.70 4.10 23.50 4.90 ;
        RECT  22.70 7.90 23.50 9.00 ;
        LAYER M1M ;
        RECT  22.75 7.85 23.45 10.55 ;
        RECT  22.85 2.75 23.55 4.95 ;
        RECT  22.65 4.05 23.55 4.95 ;
        RECT  22.65 7.85 23.55 8.90 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  25.55 2.75 26.35 4.45 ;
        RECT  25.85 2.75 26.15 10.55 ;
        RECT  25.45 7.85 26.15 10.55 ;
        RECT  25.85 2.75 26.35 8.95 ;
        RECT  25.45 7.85 26.35 8.95 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  29.65 4.10 30.55 5.00 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  36.65 5.40 37.55 6.30 ;
        END
    END J
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.25 6.65 2.55 7.35 ;
        RECT  1.65 6.65 2.55 7.65 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.30 2.50 11.00 ;
        RECT  4.05 7.95 4.75 11.00 ;
        RECT  9.80 8.20 10.50 11.00 ;
        RECT  12.30 9.55 13.00 11.00 ;
        RECT  17.15 9.05 17.85 11.00 ;
        RECT  19.85 9.15 20.55 11.00 ;
        RECT  21.40 7.90 22.10 11.00 ;
        RECT  24.10 7.90 24.80 11.00 ;
        RECT  26.80 7.90 27.50 11.00 ;
        RECT  30.35 8.50 31.05 11.00 ;
        RECT  35.20 10.65 35.90 11.00 ;
        RECT  0.00 11.00 37.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.90 2.00 1.70 3.20 ;
        RECT  4.05 2.00 4.75 4.85 ;
        RECT  2.70 2.00 5.20 2.50 ;
        RECT  8.50 2.00 9.00 4.25 ;
        RECT  9.90 3.75 10.60 4.95 ;
        RECT  8.50 3.75 13.60 4.25 ;
        RECT  12.90 3.75 13.60 5.00 ;
        RECT  18.30 2.00 18.35 5.00 ;
        RECT  17.60 4.25 18.35 5.00 ;
        RECT  18.30 2.00 18.80 4.75 ;
        RECT  17.60 4.25 18.80 4.75 ;
        RECT  19.50 2.00 20.20 2.90 ;
        RECT  21.50 2.00 22.20 4.40 ;
        RECT  24.20 2.00 24.90 4.40 ;
        RECT  26.90 2.00 27.60 4.40 ;
        RECT  29.35 2.00 30.05 3.65 ;
        RECT  34.05 2.00 34.75 3.65 ;
        RECT  0.00 0.00 37.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.25 5.35 0.75 10.25 ;
        RECT  0.25 9.55 1.15 10.25 ;
        RECT  1.00 3.80 1.80 5.85 ;
        RECT  0.25 5.35 1.80 5.85 ;
        RECT  2.70 4.20 3.55 4.90 ;
        RECT  3.05 4.20 3.55 8.85 ;
        RECT  2.70 8.15 3.55 8.85 ;
        RECT  3.05 5.55 6.35 6.05 ;
        RECT  5.35 3.20 5.85 6.05 ;
        RECT  5.85 5.55 6.35 7.40 ;
        RECT  5.85 6.70 6.55 7.40 ;
        RECT  6.40 4.20 7.55 4.90 ;
        RECT  6.85 3.00 7.55 3.70 ;
        RECT  5.35 3.20 7.55 3.70 ;
        RECT  7.05 4.20 7.55 9.25 ;
        RECT  6.40 8.55 8.00 9.25 ;
        RECT  9.35 5.65 10.05 6.35 ;
        RECT  10.35 6.90 11.05 7.60 ;
        RECT  7.05 7.10 11.05 7.60 ;
        RECT  11.40 4.75 12.10 6.15 ;
        RECT  9.35 5.65 12.10 6.15 ;
        RECT  11.60 4.75 12.10 8.85 ;
        RECT  11.15 8.10 12.10 8.85 ;
        RECT  15.25 4.30 15.50 9.85 ;
        RECT  14.80 7.15 15.50 9.85 ;
        RECT  15.25 4.30 15.75 7.65 ;
        RECT  15.25 4.30 15.95 5.00 ;
        RECT  16.95 5.95 17.65 6.70 ;
        RECT  18.50 8.15 19.20 9.85 ;
        RECT  19.00 6.95 19.70 7.65 ;
        RECT  14.80 7.15 19.70 7.65 ;
        RECT  20.00 4.35 20.70 6.45 ;
        RECT  16.95 5.95 20.70 6.45 ;
        RECT  20.20 4.35 20.70 8.65 ;
        RECT  18.50 8.15 20.70 8.65 ;
        RECT  20.00 5.75 25.35 6.25 ;
        RECT  24.65 5.55 25.35 6.25 ;
        RECT  16.95 5.95 25.35 6.25 ;
        RECT  26.80 5.25 27.50 5.95 ;
        RECT  28.25 6.45 28.95 7.20 ;
        RECT  29.35 7.50 29.85 9.25 ;
        RECT  29.00 7.65 29.85 9.25 ;
        RECT  29.35 7.50 32.40 8.00 ;
        RECT  29.00 7.65 32.40 8.00 ;
        RECT  31.70 2.95 32.40 4.80 ;
        RECT  31.70 7.50 32.40 9.15 ;
        RECT  32.60 9.65 33.30 10.35 ;
        RECT  33.05 6.45 33.75 8.15 ;
        RECT  33.40 5.25 34.10 5.95 ;
        RECT  26.80 5.45 34.10 5.95 ;
        RECT  31.70 4.30 35.10 4.80 ;
        RECT  34.40 7.50 34.90 9.15 ;
        RECT  31.70 8.65 34.90 9.15 ;
        RECT  34.60 4.30 35.10 6.95 ;
        RECT  28.25 6.45 35.10 6.95 ;
        RECT  34.40 7.50 35.10 8.25 ;
        RECT  35.40 2.95 36.10 3.65 ;
        RECT  35.60 2.95 36.10 10.15 ;
        RECT  32.60 9.65 37.25 10.15 ;
        RECT  36.55 9.65 37.25 10.35 ;
        LAYER V1M ;
        RECT  22.60 7.95 23.60 8.95 ;
        RECT  22.60 4.05 23.60 5.05 ;
    END
END JKRRX4
MACRO JKRSX1
    CLASS CORE ;
    FOREIGN JKRSX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 33.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  11.45 7.05 12.15 7.75 ;
        RECT  12.85 6.70 13.75 7.60 ;
        RECT  13.25 5.45 13.75 7.60 ;
        RECT  11.45 7.05 13.75 7.60 ;
        RECT  13.90 5.25 14.60 5.95 ;
        RECT  13.25 5.45 14.60 5.95 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M2M ;
        RECT  20.00 4.35 20.60 7.70 ;
        RECT  19.90 4.35 20.70 5.15 ;
        RECT  19.90 6.60 20.70 7.70 ;
        LAYER M1M ;
        RECT  19.95 3.75 20.65 5.20 ;
        RECT  19.95 6.70 20.65 8.90 ;
        RECT  19.85 4.30 20.75 5.20 ;
        RECT  19.85 6.70 20.75 7.60 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  22.65 3.75 23.35 4.45 ;
        RECT  22.85 3.75 23.35 8.90 ;
        RECT  22.65 6.65 23.35 8.90 ;
        RECT  22.65 6.65 23.55 7.65 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  25.45 4.10 26.35 5.00 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  32.45 5.40 33.35 6.30 ;
        END
    END J
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.25 6.65 2.55 7.35 ;
        RECT  1.65 6.65 2.55 7.65 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.30 2.50 11.00 ;
        RECT  4.05 7.95 4.75 11.00 ;
        RECT  8.75 7.90 9.45 11.00 ;
        RECT  8.00 10.45 9.60 11.00 ;
        RECT  12.05 8.70 12.75 11.00 ;
        RECT  17.05 7.40 17.75 11.00 ;
        RECT  21.30 7.10 22.00 11.00 ;
        RECT  19.20 10.45 23.50 11.00 ;
        RECT  26.15 8.50 26.85 11.00 ;
        RECT  24.90 10.10 27.40 11.00 ;
        RECT  31.00 10.65 31.70 11.00 ;
        RECT  0.00 11.00 33.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.90 2.00 1.70 3.20 ;
        RECT  4.05 2.00 4.75 4.85 ;
        RECT  8.15 2.00 9.75 3.15 ;
        RECT  9.05 2.00 9.75 4.90 ;
        RECT  11.20 2.00 11.90 3.25 ;
        RECT  17.05 2.00 17.75 3.95 ;
        RECT  21.30 2.00 22.00 4.40 ;
        RECT  25.15 2.00 25.85 3.65 ;
        RECT  29.85 2.00 30.55 3.65 ;
        RECT  0.00 0.00 33.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.25 5.35 0.75 10.25 ;
        RECT  0.25 9.55 1.20 10.25 ;
        RECT  1.00 3.80 1.80 5.85 ;
        RECT  0.25 5.35 1.80 5.85 ;
        RECT  2.70 4.20 3.55 4.90 ;
        RECT  3.05 4.20 3.55 8.85 ;
        RECT  2.70 8.15 3.55 8.85 ;
        RECT  3.05 6.70 6.55 7.20 ;
        RECT  5.35 3.20 5.85 7.20 ;
        RECT  5.85 6.70 6.55 7.40 ;
        RECT  6.40 4.20 7.55 4.90 ;
        RECT  7.05 4.20 7.10 9.55 ;
        RECT  6.40 7.90 7.10 9.55 ;
        RECT  6.85 3.00 7.55 3.70 ;
        RECT  5.35 3.20 7.55 3.70 ;
        RECT  7.05 4.20 7.55 8.40 ;
        RECT  6.40 7.90 7.55 8.40 ;
        RECT  8.30 5.45 9.00 6.15 ;
        RECT  7.05 6.70 9.95 7.20 ;
        RECT  9.25 6.70 9.95 7.40 ;
        RECT  8.30 5.45 10.95 5.95 ;
        RECT  10.45 4.35 10.95 9.45 ;
        RECT  10.45 8.75 11.25 9.45 ;
        RECT  11.55 4.15 12.25 4.85 ;
        RECT  10.45 4.35 12.25 4.85 ;
        RECT  13.70 3.30 14.40 4.00 ;
        RECT  13.70 3.45 15.60 4.00 ;
        RECT  14.55 7.20 15.10 10.50 ;
        RECT  14.40 8.70 15.10 10.50 ;
        RECT  15.10 3.45 15.60 7.90 ;
        RECT  14.55 7.20 15.60 7.90 ;
        RECT  16.60 4.45 17.30 5.15 ;
        RECT  17.40 5.70 18.10 6.40 ;
        RECT  15.10 5.90 18.10 6.40 ;
        RECT  18.40 3.25 19.10 4.95 ;
        RECT  16.60 4.45 19.10 4.95 ;
        RECT  18.40 7.40 19.15 8.15 ;
        RECT  18.65 3.25 19.10 9.95 ;
        RECT  18.60 3.25 19.10 8.15 ;
        RECT  18.65 5.70 19.15 9.95 ;
        RECT  18.65 9.25 19.35 9.95 ;
        RECT  21.65 5.50 22.35 6.20 ;
        RECT  18.60 5.70 22.35 6.20 ;
        RECT  24.05 5.25 24.75 6.00 ;
        RECT  24.05 6.50 24.75 7.25 ;
        RECT  25.15 7.50 25.65 9.20 ;
        RECT  24.80 8.50 25.65 9.20 ;
        RECT  25.15 7.50 28.20 8.00 ;
        RECT  27.50 2.95 28.20 4.65 ;
        RECT  27.50 7.50 28.20 9.15 ;
        RECT  28.40 9.65 29.10 10.35 ;
        RECT  28.85 6.50 29.55 8.15 ;
        RECT  29.20 5.30 29.90 6.00 ;
        RECT  24.05 5.50 29.90 6.00 ;
        RECT  27.50 4.15 30.85 4.65 ;
        RECT  30.20 7.50 30.70 9.15 ;
        RECT  27.50 8.65 30.70 9.15 ;
        RECT  30.35 4.15 30.85 7.00 ;
        RECT  24.05 6.50 30.85 7.00 ;
        RECT  30.20 7.50 30.90 8.25 ;
        RECT  31.20 2.95 31.90 3.65 ;
        RECT  31.40 2.95 31.90 10.15 ;
        RECT  28.40 9.65 33.05 10.15 ;
        RECT  32.35 9.65 33.05 10.35 ;
        LAYER V1M ;
        RECT  19.80 6.65 20.80 7.65 ;
        RECT  19.80 4.05 20.80 5.05 ;
    END
END JKRSX1
MACRO JKRSX2
    CLASS CORE ;
    FOREIGN JKRSX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 33.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  11.45 7.05 12.15 7.75 ;
        RECT  12.85 6.70 13.75 7.60 ;
        RECT  13.25 5.45 13.75 7.60 ;
        RECT  11.45 7.05 13.75 7.60 ;
        RECT  13.90 5.25 14.60 5.95 ;
        RECT  13.25 5.45 14.60 5.95 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M2M ;
        RECT  20.00 4.35 20.60 7.70 ;
        RECT  19.90 4.35 20.70 5.15 ;
        RECT  19.90 6.60 20.70 7.70 ;
        LAYER M1M ;
        RECT  19.95 2.70 20.65 5.20 ;
        RECT  19.95 6.70 20.65 10.55 ;
        RECT  19.85 4.30 20.75 5.20 ;
        RECT  19.85 6.70 20.75 7.60 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  22.65 2.70 23.35 4.45 ;
        RECT  22.85 2.70 23.35 10.55 ;
        RECT  22.65 6.65 23.35 10.55 ;
        RECT  22.65 6.65 23.55 7.65 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  25.45 4.10 26.35 5.00 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  32.45 5.40 33.35 6.30 ;
        END
    END J
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.25 6.65 2.55 7.35 ;
        RECT  1.65 6.65 2.55 7.65 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.30 2.50 11.00 ;
        RECT  4.05 7.95 4.75 11.00 ;
        RECT  8.75 7.90 9.45 11.00 ;
        RECT  8.00 10.45 9.60 11.00 ;
        RECT  12.05 8.70 12.75 11.00 ;
        RECT  17.05 7.40 17.75 11.00 ;
        RECT  21.30 7.25 22.00 11.00 ;
        RECT  26.15 8.50 26.85 11.00 ;
        RECT  24.90 10.10 27.40 11.00 ;
        RECT  31.00 10.65 31.70 11.00 ;
        RECT  0.00 11.00 33.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.90 2.00 1.70 3.20 ;
        RECT  4.05 2.00 4.75 4.85 ;
        RECT  8.15 2.00 9.75 3.15 ;
        RECT  9.05 2.00 9.75 4.90 ;
        RECT  11.20 2.00 11.90 3.25 ;
        RECT  17.05 2.00 17.75 3.95 ;
        RECT  21.30 2.00 22.00 4.40 ;
        RECT  25.15 2.00 25.85 3.65 ;
        RECT  29.85 2.00 30.55 3.65 ;
        RECT  0.00 0.00 33.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.25 5.35 0.75 10.25 ;
        RECT  0.25 9.55 1.20 10.25 ;
        RECT  1.00 3.80 1.80 5.85 ;
        RECT  0.25 5.35 1.80 5.85 ;
        RECT  2.70 4.20 3.55 4.90 ;
        RECT  3.05 4.20 3.55 8.85 ;
        RECT  2.70 8.15 3.55 8.85 ;
        RECT  3.05 6.70 6.55 7.20 ;
        RECT  5.35 3.20 5.85 7.20 ;
        RECT  5.85 6.70 6.55 7.40 ;
        RECT  6.40 4.20 7.55 4.90 ;
        RECT  7.05 4.20 7.10 9.55 ;
        RECT  6.40 7.90 7.10 9.55 ;
        RECT  6.85 3.00 7.55 3.70 ;
        RECT  5.35 3.20 7.55 3.70 ;
        RECT  7.05 4.20 7.55 8.40 ;
        RECT  6.40 7.90 7.55 8.40 ;
        RECT  8.30 5.45 9.00 6.15 ;
        RECT  7.05 6.70 9.95 7.20 ;
        RECT  9.25 6.70 9.95 7.40 ;
        RECT  8.30 5.45 10.95 5.95 ;
        RECT  10.45 4.35 10.95 9.45 ;
        RECT  10.45 8.75 11.25 9.45 ;
        RECT  11.55 4.15 12.25 4.85 ;
        RECT  10.45 4.35 12.25 4.85 ;
        RECT  13.70 3.30 14.40 4.00 ;
        RECT  13.70 3.45 15.60 4.00 ;
        RECT  14.55 7.20 15.10 10.50 ;
        RECT  14.40 8.70 15.10 10.50 ;
        RECT  15.10 3.45 15.60 7.90 ;
        RECT  14.55 7.20 15.60 7.90 ;
        RECT  16.60 4.45 17.30 5.15 ;
        RECT  17.40 5.70 18.10 6.40 ;
        RECT  15.10 5.90 18.10 6.40 ;
        RECT  18.40 3.25 19.10 4.95 ;
        RECT  16.60 4.45 19.10 4.95 ;
        RECT  18.40 7.40 19.15 8.15 ;
        RECT  18.65 3.25 19.10 9.95 ;
        RECT  18.60 3.25 19.10 8.15 ;
        RECT  18.65 5.70 19.15 9.95 ;
        RECT  18.65 9.25 19.35 9.95 ;
        RECT  21.65 5.50 22.35 6.20 ;
        RECT  18.60 5.70 22.35 6.20 ;
        RECT  24.05 5.25 24.75 6.00 ;
        RECT  24.05 6.50 24.75 7.25 ;
        RECT  25.15 7.50 25.65 9.20 ;
        RECT  24.80 8.50 25.65 9.20 ;
        RECT  25.15 7.50 28.20 8.00 ;
        RECT  27.50 2.95 28.20 4.65 ;
        RECT  27.50 7.50 28.20 9.15 ;
        RECT  28.40 9.65 29.10 10.35 ;
        RECT  28.85 6.50 29.55 8.15 ;
        RECT  29.20 5.30 29.90 6.00 ;
        RECT  24.05 5.50 29.90 6.00 ;
        RECT  27.50 4.15 30.85 4.65 ;
        RECT  30.20 7.50 30.70 9.15 ;
        RECT  27.50 8.65 30.70 9.15 ;
        RECT  30.35 4.15 30.85 7.00 ;
        RECT  24.05 6.50 30.85 7.00 ;
        RECT  30.20 7.50 30.90 8.25 ;
        RECT  31.20 2.95 31.90 3.65 ;
        RECT  31.40 2.95 31.90 10.15 ;
        RECT  28.40 9.65 33.05 10.15 ;
        RECT  32.35 9.65 33.05 10.35 ;
        LAYER V1M ;
        RECT  19.80 6.65 20.80 7.65 ;
        RECT  19.80 4.05 20.80 5.05 ;
    END
END JKRSX2
MACRO JKRSX4
    CLASS CORE ;
    FOREIGN JKRSX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 36.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  11.45 7.05 12.15 7.75 ;
        RECT  12.85 6.70 13.75 7.60 ;
        RECT  13.25 5.45 13.75 7.60 ;
        RECT  11.45 7.05 13.75 7.60 ;
        RECT  13.90 5.25 14.60 5.95 ;
        RECT  13.25 5.45 14.60 5.95 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M2M ;
        RECT  21.40 4.35 22.00 7.70 ;
        RECT  21.30 4.35 22.10 5.15 ;
        RECT  21.30 6.60 22.10 7.70 ;
        LAYER M1M ;
        RECT  21.35 2.70 22.05 5.20 ;
        RECT  21.35 6.70 22.05 10.55 ;
        RECT  21.25 4.30 22.15 5.20 ;
        RECT  21.25 6.70 22.15 7.60 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  24.05 2.70 24.75 4.45 ;
        RECT  24.25 2.70 24.75 10.55 ;
        RECT  24.05 6.65 24.75 10.55 ;
        RECT  24.05 6.65 24.95 7.65 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  28.25 4.10 29.15 5.00 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  35.25 5.40 36.15 6.30 ;
        END
    END J
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.25 6.65 2.55 7.35 ;
        RECT  1.65 6.65 2.55 7.65 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.30 2.50 11.00 ;
        RECT  4.05 7.95 4.75 11.00 ;
        RECT  8.75 7.90 9.45 11.00 ;
        RECT  8.00 10.45 9.60 11.00 ;
        RECT  12.05 8.70 12.75 11.00 ;
        RECT  17.05 7.40 17.75 11.00 ;
        RECT  20.00 7.25 20.70 11.00 ;
        RECT  22.70 7.25 23.40 11.00 ;
        RECT  25.40 7.25 26.10 11.00 ;
        RECT  28.95 8.50 29.65 11.00 ;
        RECT  27.70 10.10 30.20 11.00 ;
        RECT  33.80 10.65 34.50 11.00 ;
        RECT  0.00 11.00 36.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.90 2.00 1.70 3.20 ;
        RECT  4.05 2.00 4.75 4.85 ;
        RECT  8.15 2.00 9.75 3.15 ;
        RECT  9.05 2.00 9.75 4.90 ;
        RECT  11.20 2.00 11.90 3.25 ;
        RECT  17.05 2.00 17.75 3.95 ;
        RECT  20.00 2.00 20.70 4.40 ;
        RECT  22.70 2.00 23.40 4.40 ;
        RECT  25.40 2.00 26.10 4.40 ;
        RECT  27.95 2.00 28.65 3.65 ;
        RECT  32.65 2.00 33.35 3.65 ;
        RECT  0.00 0.00 36.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.25 5.35 0.75 10.25 ;
        RECT  0.25 9.55 1.20 10.25 ;
        RECT  1.00 3.80 1.80 5.85 ;
        RECT  0.25 5.35 1.80 5.85 ;
        RECT  2.70 4.20 3.55 4.90 ;
        RECT  3.05 4.20 3.55 8.85 ;
        RECT  2.70 8.15 3.55 8.85 ;
        RECT  3.05 6.70 6.55 7.20 ;
        RECT  5.35 3.20 5.85 7.20 ;
        RECT  5.85 6.70 6.55 7.40 ;
        RECT  6.40 4.20 7.55 4.90 ;
        RECT  7.05 4.20 7.10 9.55 ;
        RECT  6.40 7.90 7.10 9.55 ;
        RECT  6.85 3.00 7.55 3.70 ;
        RECT  5.35 3.20 7.55 3.70 ;
        RECT  7.05 4.20 7.55 8.40 ;
        RECT  6.40 7.90 7.55 8.40 ;
        RECT  8.30 5.45 9.00 6.15 ;
        RECT  7.05 6.70 9.95 7.20 ;
        RECT  9.25 6.70 9.95 7.40 ;
        RECT  8.30 5.45 10.95 5.95 ;
        RECT  10.45 4.35 10.95 9.45 ;
        RECT  10.45 8.75 11.25 9.45 ;
        RECT  11.55 4.15 12.25 4.85 ;
        RECT  10.45 4.35 12.25 4.85 ;
        RECT  13.70 3.30 14.40 4.00 ;
        RECT  13.70 3.45 15.60 4.00 ;
        RECT  14.55 7.20 15.10 10.50 ;
        RECT  14.40 8.70 15.10 10.50 ;
        RECT  15.10 3.45 15.60 7.90 ;
        RECT  14.55 7.20 15.60 7.90 ;
        RECT  16.60 4.45 17.30 5.15 ;
        RECT  17.40 5.70 18.10 6.40 ;
        RECT  15.10 5.90 18.10 6.40 ;
        RECT  18.40 3.25 19.10 4.95 ;
        RECT  16.60 4.45 19.10 4.95 ;
        RECT  18.40 7.40 19.15 8.15 ;
        RECT  18.65 3.25 19.10 9.95 ;
        RECT  18.60 3.25 19.10 8.15 ;
        RECT  18.65 5.70 19.15 9.95 ;
        RECT  18.65 9.25 19.35 9.95 ;
        RECT  23.05 5.50 23.75 6.20 ;
        RECT  18.60 5.70 23.75 6.20 ;
        RECT  26.85 5.25 27.55 6.00 ;
        RECT  26.85 6.50 27.55 7.25 ;
        RECT  27.95 7.50 28.45 9.20 ;
        RECT  27.60 8.50 28.45 9.20 ;
        RECT  27.95 7.50 31.00 8.00 ;
        RECT  30.30 2.95 31.00 4.65 ;
        RECT  30.30 7.50 31.00 9.15 ;
        RECT  31.20 9.65 31.90 10.35 ;
        RECT  31.65 6.50 32.35 8.15 ;
        RECT  32.00 5.30 32.70 6.00 ;
        RECT  26.85 5.50 32.70 6.00 ;
        RECT  30.30 4.15 33.65 4.65 ;
        RECT  33.00 7.50 33.50 9.15 ;
        RECT  30.30 8.65 33.50 9.15 ;
        RECT  33.15 4.15 33.65 7.00 ;
        RECT  26.85 6.50 33.65 7.00 ;
        RECT  33.00 7.50 33.70 8.25 ;
        RECT  34.00 2.95 34.70 3.65 ;
        RECT  34.20 2.95 34.70 10.15 ;
        RECT  31.20 9.65 35.85 10.15 ;
        RECT  35.15 9.65 35.85 10.35 ;
        LAYER V1M ;
        RECT  21.20 6.65 22.20 7.65 ;
        RECT  21.20 4.05 22.20 5.05 ;
    END
END JKRSX4
MACRO LGCNX1
    CLASS CORE ;
    FOREIGN LGCNX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  15.50 3.75 16.35 4.45 ;
        RECT  15.85 3.75 16.35 8.90 ;
        RECT  15.65 7.10 16.35 8.90 ;
        RECT  15.65 8.00 16.55 8.90 ;
        END
    END GCLK
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 4.10 6.75 5.00 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.80 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END CLK
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.45 2.50 11.00 ;
        RECT  6.65 6.55 7.35 11.00 ;
        RECT  6.50 8.35 7.35 11.00 ;
        RECT  4.95 10.75 8.05 11.00 ;
        RECT  10.30 9.00 11.00 11.00 ;
        RECT  14.15 7.10 14.85 11.00 ;
        RECT  15.65 10.10 16.35 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.95 2.00 2.65 4.50 ;
        RECT  1.80 3.80 2.65 4.50 ;
        RECT  6.65 2.00 7.20 3.65 ;
        RECT  6.65 2.95 7.35 3.65 ;
        RECT  11.30 2.00 12.00 4.50 ;
        RECT  11.30 3.80 12.15 4.50 ;
        RECT  14.15 2.00 14.85 4.45 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.80 0.95 9.05 ;
        RECT  0.45 3.80 1.15 4.50 ;
        RECT  0.45 7.45 1.15 9.05 ;
        RECT  1.40 6.20 2.10 6.90 ;
        RECT  2.25 4.95 2.95 5.65 ;
        RECT  0.45 5.15 2.95 5.65 ;
        RECT  1.40 6.40 4.65 6.90 ;
        RECT  3.80 4.30 4.30 6.90 ;
        RECT  4.15 6.40 4.65 9.00 ;
        RECT  4.30 3.00 4.80 4.80 ;
        RECT  3.80 4.30 4.80 4.80 ;
        RECT  4.15 7.40 4.85 9.00 ;
        RECT  4.30 3.00 5.00 3.70 ;
        RECT  4.75 5.25 5.45 5.95 ;
        RECT  4.75 5.45 8.40 5.95 ;
        RECT  7.90 3.00 8.40 8.10 ;
        RECT  7.90 3.00 8.70 3.70 ;
        RECT  7.90 6.50 8.70 8.10 ;
        RECT  8.85 4.15 9.65 4.85 ;
        RECT  9.15 3.00 9.65 10.55 ;
        RECT  8.95 8.95 9.65 10.55 ;
        RECT  9.15 3.00 10.65 3.70 ;
        RECT  11.80 7.10 12.50 10.55 ;
        RECT  12.80 3.75 13.50 4.45 ;
        RECT  13.00 3.75 13.50 7.60 ;
        RECT  11.80 7.10 13.50 7.60 ;
        RECT  13.00 5.45 15.40 5.95 ;
        RECT  14.70 5.45 15.40 6.15 ;
    END
END LGCNX1
MACRO LGCNX2
    CLASS CORE ;
    FOREIGN LGCNX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  15.65 2.75 16.35 4.45 ;
        RECT  15.85 2.75 16.35 10.55 ;
        RECT  15.65 7.10 16.35 10.55 ;
        RECT  15.65 8.00 16.55 8.90 ;
        END
    END GCLK
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 4.10 6.75 5.00 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.80 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END CLK
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.45 2.50 11.00 ;
        RECT  6.65 6.55 7.35 11.00 ;
        RECT  6.50 8.35 7.35 11.00 ;
        RECT  4.85 10.75 8.25 11.00 ;
        RECT  10.45 9.00 11.15 11.00 ;
        RECT  14.30 7.10 15.00 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.95 2.00 2.65 4.50 ;
        RECT  1.80 3.80 2.65 4.50 ;
        RECT  6.65 2.00 7.35 3.65 ;
        RECT  11.30 2.00 12.00 4.50 ;
        RECT  11.30 3.80 12.15 4.50 ;
        RECT  14.30 2.00 15.00 4.45 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.80 0.95 9.05 ;
        RECT  0.45 3.80 1.15 4.50 ;
        RECT  0.45 7.45 1.15 9.05 ;
        RECT  1.40 6.20 2.10 6.90 ;
        RECT  2.25 4.95 2.95 5.65 ;
        RECT  0.45 5.15 2.95 5.65 ;
        RECT  1.40 6.40 4.65 6.90 ;
        RECT  3.80 4.30 4.30 6.90 ;
        RECT  4.15 6.40 4.65 9.00 ;
        RECT  4.30 3.00 4.80 4.80 ;
        RECT  3.80 4.30 4.80 4.80 ;
        RECT  4.15 7.40 4.85 9.00 ;
        RECT  4.30 3.00 5.00 3.70 ;
        RECT  4.75 5.25 5.45 5.95 ;
        RECT  4.75 5.45 8.40 5.95 ;
        RECT  7.90 3.00 8.40 8.10 ;
        RECT  7.90 3.00 8.70 3.70 ;
        RECT  7.90 6.50 8.70 8.10 ;
        RECT  8.85 4.15 9.80 4.85 ;
        RECT  9.30 3.00 9.80 10.55 ;
        RECT  9.10 8.95 9.80 10.55 ;
        RECT  9.30 3.00 10.65 3.70 ;
        RECT  11.95 7.10 12.65 10.55 ;
        RECT  12.80 3.75 13.50 4.45 ;
        RECT  13.00 3.75 13.50 7.60 ;
        RECT  11.95 7.10 13.50 7.60 ;
        RECT  13.00 5.25 15.40 5.75 ;
        RECT  14.70 5.25 15.40 5.95 ;
    END
END LGCNX2
MACRO LGCNX3
    CLASS CORE ;
    FOREIGN LGCNX3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  15.50 3.50 16.35 4.20 ;
        RECT  15.85 3.50 16.35 9.85 ;
        RECT  15.65 7.10 16.35 9.85 ;
        RECT  15.65 8.00 16.55 8.90 ;
        END
    END GCLK
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 4.10 6.75 5.00 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.80 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END CLK
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.45 2.50 11.00 ;
        RECT  6.65 6.55 7.35 11.00 ;
        RECT  6.50 8.35 7.35 11.00 ;
        RECT  4.95 10.75 8.05 11.00 ;
        RECT  10.30 9.00 11.00 11.00 ;
        RECT  14.15 7.10 14.85 11.00 ;
        RECT  17.00 7.10 17.70 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.95 2.00 2.65 4.50 ;
        RECT  1.80 3.80 2.65 4.50 ;
        RECT  6.65 2.00 7.20 3.65 ;
        RECT  6.65 2.95 7.35 3.65 ;
        RECT  11.30 2.00 12.00 4.50 ;
        RECT  11.30 3.80 12.15 4.50 ;
        RECT  14.15 2.00 14.85 4.45 ;
        RECT  16.85 2.00 17.55 4.45 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.80 0.95 9.05 ;
        RECT  0.45 3.80 1.15 4.50 ;
        RECT  0.45 7.45 1.15 9.05 ;
        RECT  1.40 6.20 2.10 6.90 ;
        RECT  2.25 4.95 2.95 5.65 ;
        RECT  0.45 5.15 2.95 5.65 ;
        RECT  1.40 6.40 4.65 6.90 ;
        RECT  3.80 4.30 4.30 6.90 ;
        RECT  4.15 6.40 4.65 9.00 ;
        RECT  4.30 3.00 4.80 4.80 ;
        RECT  3.80 4.30 4.80 4.80 ;
        RECT  4.15 7.40 4.85 9.00 ;
        RECT  4.30 3.00 5.00 3.70 ;
        RECT  4.75 5.25 5.45 5.95 ;
        RECT  4.75 5.45 8.40 5.95 ;
        RECT  7.90 3.00 8.40 8.10 ;
        RECT  7.90 3.00 8.70 3.70 ;
        RECT  7.90 6.50 8.70 8.10 ;
        RECT  8.85 4.15 9.65 4.85 ;
        RECT  9.15 3.00 9.65 10.55 ;
        RECT  8.95 8.95 9.65 10.55 ;
        RECT  9.15 3.00 10.65 3.70 ;
        RECT  11.80 7.10 12.50 10.55 ;
        RECT  12.80 3.75 13.50 4.45 ;
        RECT  13.00 3.75 13.50 7.60 ;
        RECT  11.80 7.10 13.50 7.60 ;
        RECT  13.00 5.45 15.40 5.95 ;
        RECT  14.70 5.45 15.40 6.15 ;
    END
END LGCNX3
MACRO LGCNX4
    CLASS CORE ;
    FOREIGN LGCNX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  15.65 2.75 16.35 4.45 ;
        RECT  15.85 2.75 16.35 10.55 ;
        RECT  15.65 7.10 16.35 10.55 ;
        RECT  15.65 8.00 16.55 8.90 ;
        END
    END GCLK
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 4.10 6.75 5.00 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.80 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END CLK
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.45 2.50 11.00 ;
        RECT  6.65 6.55 7.35 11.00 ;
        RECT  6.50 8.35 7.35 11.00 ;
        RECT  4.85 10.75 8.25 11.00 ;
        RECT  10.45 9.00 11.15 11.00 ;
        RECT  14.30 7.10 15.00 11.00 ;
        RECT  17.00 7.10 17.70 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.95 2.00 2.65 4.50 ;
        RECT  1.80 3.80 2.65 4.50 ;
        RECT  6.65 2.00 7.35 3.65 ;
        RECT  11.30 2.00 12.00 4.50 ;
        RECT  11.30 3.80 12.15 4.50 ;
        RECT  14.30 2.00 15.00 4.45 ;
        RECT  17.00 2.00 17.70 4.45 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.80 0.95 9.05 ;
        RECT  0.45 3.80 1.15 4.50 ;
        RECT  0.45 7.45 1.15 9.05 ;
        RECT  1.40 6.20 2.10 6.90 ;
        RECT  2.25 4.95 2.95 5.65 ;
        RECT  0.45 5.15 2.95 5.65 ;
        RECT  1.40 6.40 4.65 6.90 ;
        RECT  3.80 4.30 4.30 6.90 ;
        RECT  4.15 6.40 4.65 9.00 ;
        RECT  4.30 3.00 4.80 4.80 ;
        RECT  3.80 4.30 4.80 4.80 ;
        RECT  4.15 7.40 4.85 9.00 ;
        RECT  4.30 3.00 5.00 3.70 ;
        RECT  4.75 5.25 5.45 5.95 ;
        RECT  4.75 5.45 8.40 5.95 ;
        RECT  7.90 3.00 8.40 8.10 ;
        RECT  7.90 3.00 8.70 3.70 ;
        RECT  7.90 6.50 8.70 8.10 ;
        RECT  8.85 4.15 9.80 4.85 ;
        RECT  9.30 3.00 9.80 10.55 ;
        RECT  9.10 8.95 9.80 10.55 ;
        RECT  9.30 3.00 10.65 3.70 ;
        RECT  11.95 7.10 12.65 10.55 ;
        RECT  12.80 3.75 13.50 4.45 ;
        RECT  13.00 3.75 13.50 7.60 ;
        RECT  11.95 7.10 13.50 7.60 ;
        RECT  13.00 5.25 15.40 5.75 ;
        RECT  14.70 5.25 15.40 5.95 ;
    END
END LGCNX4
MACRO LGCNX8
    CLASS CORE ;
    FOREIGN LGCNX8 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  18.55 2.75 19.25 4.45 ;
        RECT  18.75 2.75 19.25 10.55 ;
        RECT  18.55 7.10 19.25 10.55 ;
        RECT  19.85 5.40 20.75 6.30 ;
        RECT  18.75 5.40 21.75 5.90 ;
        RECT  21.25 2.75 21.75 10.55 ;
        RECT  21.25 2.75 21.95 4.45 ;
        RECT  21.25 7.10 21.95 10.55 ;
        END
    END GCLK
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 4.10 6.75 5.00 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.55 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.35 12.35 6.30 ;
        END
    END CLK
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.45 2.50 11.00 ;
        RECT  6.65 6.45 7.35 11.00 ;
        RECT  6.50 8.30 7.35 11.00 ;
        RECT  10.15 9.00 10.85 11.00 ;
        RECT  14.00 7.10 17.90 7.80 ;
        RECT  17.20 7.10 17.90 11.00 ;
        RECT  19.90 7.10 20.60 11.00 ;
        RECT  22.60 7.10 23.30 11.00 ;
        RECT  0.00 11.00 23.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.95 2.00 2.65 4.50 ;
        RECT  1.80 3.80 2.65 4.50 ;
        RECT  6.65 2.00 7.35 3.65 ;
        RECT  11.65 2.00 12.35 3.65 ;
        RECT  14.35 2.00 15.05 3.65 ;
        RECT  17.20 2.00 17.90 4.45 ;
        RECT  19.90 2.00 20.60 4.45 ;
        RECT  22.60 2.00 23.30 4.45 ;
        RECT  0.00 0.00 23.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.80 0.95 9.05 ;
        RECT  0.45 3.80 1.15 4.50 ;
        RECT  0.45 7.45 1.15 9.05 ;
        RECT  1.40 6.20 2.10 6.90 ;
        RECT  2.25 4.95 2.95 5.65 ;
        RECT  0.45 5.15 2.95 5.65 ;
        RECT  1.40 6.40 4.65 6.90 ;
        RECT  3.80 4.30 4.30 6.90 ;
        RECT  4.15 6.40 4.65 9.00 ;
        RECT  4.30 3.00 4.80 4.80 ;
        RECT  3.80 4.30 4.80 4.80 ;
        RECT  4.15 7.40 4.85 9.00 ;
        RECT  4.30 3.00 5.00 3.70 ;
        RECT  4.75 5.25 5.45 5.95 ;
        RECT  4.75 5.45 8.40 5.95 ;
        RECT  7.90 3.00 8.40 8.00 ;
        RECT  7.90 3.00 8.70 3.70 ;
        RECT  7.90 6.40 8.70 8.00 ;
        RECT  8.85 4.15 9.65 4.85 ;
        RECT  9.15 2.95 9.65 10.55 ;
        RECT  8.80 8.95 9.65 10.55 ;
        RECT  9.15 2.95 11.00 3.65 ;
        RECT  11.65 7.10 12.35 10.15 ;
        RECT  13.00 2.95 13.50 7.60 ;
        RECT  11.65 7.10 13.50 7.60 ;
        RECT  13.00 2.95 13.70 3.65 ;
        RECT  11.65 9.45 15.55 10.15 ;
        RECT  15.70 2.95 16.20 5.75 ;
        RECT  15.70 2.95 16.40 3.65 ;
        RECT  13.00 5.25 18.30 5.75 ;
        RECT  17.60 5.25 18.30 5.95 ;
    END
END LGCNX8
MACRO LGCPX1
    CLASS CORE ;
    FOREIGN LGCPX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  14.25 3.75 14.95 4.45 ;
        RECT  14.45 3.75 14.95 9.10 ;
        RECT  14.25 7.30 14.95 9.10 ;
        RECT  14.25 8.00 15.15 9.10 ;
        END
    END GCLK
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END CLK
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.70 2.50 11.00 ;
        RECT  0.45 10.25 2.50 11.00 ;
        RECT  6.50 7.70 7.20 11.00 ;
        RECT  10.05 7.30 10.75 9.25 ;
        RECT  10.05 8.55 12.00 9.25 ;
        RECT  11.30 8.55 12.00 11.00 ;
        RECT  12.90 7.30 13.60 11.00 ;
        RECT  12.90 10.10 14.95 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.50 ;
        RECT  6.50 2.00 7.20 4.65 ;
        RECT  12.90 2.00 13.60 4.50 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.65 7.70 4.85 8.20 ;
        RECT  0.45 3.80 0.95 9.30 ;
        RECT  0.45 3.80 1.15 4.50 ;
        RECT  0.45 7.70 1.15 9.30 ;
        RECT  1.40 6.45 2.10 7.15 ;
        RECT  2.25 4.95 2.95 5.65 ;
        RECT  0.45 5.15 2.95 5.65 ;
        RECT  1.40 6.65 4.15 7.15 ;
        RECT  3.65 3.85 4.15 8.20 ;
        RECT  3.65 3.85 4.85 4.55 ;
        RECT  4.15 7.70 4.85 9.30 ;
        RECT  4.60 6.25 5.30 7.25 ;
        RECT  4.60 6.75 8.35 7.25 ;
        RECT  7.85 3.95 8.35 9.10 ;
        RECT  7.85 3.95 8.55 4.65 ;
        RECT  7.85 7.50 8.55 9.10 ;
        RECT  8.90 2.45 9.60 3.15 ;
        RECT  8.80 5.45 9.60 6.15 ;
        RECT  9.10 2.45 9.60 10.55 ;
        RECT  8.95 9.85 10.60 10.55 ;
        RECT  10.55 3.75 11.25 4.45 ;
        RECT  10.55 3.95 12.10 4.45 ;
        RECT  11.60 3.95 12.10 8.00 ;
        RECT  11.40 7.30 12.10 8.00 ;
        RECT  11.60 5.65 14.00 6.15 ;
        RECT  13.30 5.65 14.00 6.35 ;
    END
END LGCPX1
MACRO LGCPX2
    CLASS CORE ;
    FOREIGN LGCPX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  14.25 2.75 14.95 4.45 ;
        RECT  14.45 2.75 14.95 10.55 ;
        RECT  14.25 7.15 14.95 10.55 ;
        RECT  14.25 8.00 15.15 9.10 ;
        END
    END GCLK
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END CLK
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.70 2.50 11.00 ;
        RECT  0.45 10.25 2.50 11.00 ;
        RECT  6.50 7.70 7.20 11.00 ;
        RECT  10.05 7.30 10.75 9.25 ;
        RECT  10.05 8.55 12.00 9.25 ;
        RECT  11.30 8.55 12.00 11.00 ;
        RECT  12.90 7.30 13.60 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.50 ;
        RECT  6.50 2.00 7.20 4.65 ;
        RECT  12.90 2.00 13.60 4.45 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.65 7.70 4.85 8.20 ;
        RECT  0.45 3.80 0.95 9.30 ;
        RECT  0.45 3.80 1.15 4.50 ;
        RECT  0.45 7.70 1.15 9.30 ;
        RECT  1.40 6.45 2.10 7.15 ;
        RECT  2.25 4.95 2.95 5.65 ;
        RECT  0.45 5.15 2.95 5.65 ;
        RECT  1.40 6.65 4.15 7.15 ;
        RECT  3.65 3.85 4.15 8.20 ;
        RECT  3.65 3.85 4.85 4.55 ;
        RECT  4.15 7.70 4.85 9.30 ;
        RECT  4.60 6.25 5.30 7.25 ;
        RECT  4.60 6.75 8.35 7.25 ;
        RECT  7.85 3.95 8.35 9.10 ;
        RECT  7.85 3.95 8.55 4.65 ;
        RECT  7.85 7.50 8.55 9.10 ;
        RECT  8.90 2.45 9.60 3.15 ;
        RECT  8.80 5.45 9.60 6.15 ;
        RECT  9.10 2.45 9.60 10.55 ;
        RECT  8.95 9.85 10.60 10.55 ;
        RECT  10.40 3.75 11.10 4.45 ;
        RECT  10.40 3.95 12.10 4.45 ;
        RECT  11.60 3.95 12.10 8.00 ;
        RECT  11.40 7.30 12.10 8.00 ;
        RECT  11.60 5.65 14.00 6.15 ;
        RECT  13.30 5.65 14.00 6.35 ;
    END
END LGCPX2
MACRO LGCPX3
    CLASS CORE ;
    FOREIGN LGCPX3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  14.25 3.50 14.95 4.20 ;
        RECT  14.45 3.50 14.95 9.65 ;
        RECT  14.25 7.15 14.95 9.65 ;
        RECT  14.25 8.00 15.15 9.10 ;
        END
    END GCLK
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END CLK
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.70 2.50 11.00 ;
        RECT  0.45 10.25 2.50 11.00 ;
        RECT  6.50 7.70 7.20 11.00 ;
        RECT  10.05 7.30 10.75 9.40 ;
        RECT  10.05 8.70 12.00 9.40 ;
        RECT  11.30 8.70 12.00 11.00 ;
        RECT  12.90 7.30 13.60 11.00 ;
        RECT  15.60 7.30 16.30 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.50 ;
        RECT  6.50 2.00 7.20 4.65 ;
        RECT  12.75 2.00 13.45 4.45 ;
        RECT  15.60 2.00 16.30 4.20 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.65 7.70 4.85 8.20 ;
        RECT  0.45 3.80 0.95 9.30 ;
        RECT  0.45 3.80 1.15 4.50 ;
        RECT  0.45 7.70 1.15 9.30 ;
        RECT  1.40 6.45 2.10 7.15 ;
        RECT  2.25 4.95 2.95 5.65 ;
        RECT  0.45 5.15 2.95 5.65 ;
        RECT  1.40 6.65 4.15 7.15 ;
        RECT  3.65 3.85 4.15 8.20 ;
        RECT  3.65 3.85 4.85 4.55 ;
        RECT  4.15 7.70 4.85 9.30 ;
        RECT  4.60 6.25 5.30 7.25 ;
        RECT  4.60 6.75 8.35 7.25 ;
        RECT  7.85 3.95 8.35 9.10 ;
        RECT  7.85 3.95 8.55 4.65 ;
        RECT  7.85 7.50 8.55 9.10 ;
        RECT  8.85 2.45 9.55 3.15 ;
        RECT  8.80 5.45 9.55 6.15 ;
        RECT  9.05 2.45 9.55 10.55 ;
        RECT  8.95 9.85 10.60 10.55 ;
        RECT  10.40 2.75 11.10 4.45 ;
        RECT  10.40 3.95 12.10 4.45 ;
        RECT  11.60 3.95 12.10 8.25 ;
        RECT  11.40 7.55 12.10 8.25 ;
        RECT  11.60 5.65 14.00 6.15 ;
        RECT  13.30 5.65 14.00 6.35 ;
    END
END LGCPX3
MACRO LGCPX4
    CLASS CORE ;
    FOREIGN LGCPX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  14.10 2.75 14.80 4.45 ;
        RECT  14.30 2.75 14.80 10.55 ;
        RECT  14.25 7.15 14.95 10.55 ;
        RECT  14.25 8.00 15.15 8.90 ;
        END
    END GCLK
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END CLK
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.70 2.50 11.00 ;
        RECT  0.45 10.30 2.50 11.00 ;
        RECT  6.50 7.70 7.20 11.00 ;
        RECT  10.05 7.30 10.75 9.40 ;
        RECT  10.05 8.70 12.00 9.40 ;
        RECT  11.30 8.70 12.00 11.00 ;
        RECT  12.90 7.30 13.60 11.00 ;
        RECT  15.60 7.30 16.30 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.50 ;
        RECT  6.50 2.00 7.20 4.65 ;
        RECT  12.75 2.00 13.45 4.45 ;
        RECT  15.45 2.00 16.15 4.45 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.65 7.70 4.85 8.20 ;
        RECT  0.45 3.80 0.95 9.30 ;
        RECT  0.45 3.80 1.15 4.50 ;
        RECT  0.45 7.70 1.15 9.30 ;
        RECT  1.40 6.45 2.10 7.15 ;
        RECT  2.25 4.95 2.95 5.65 ;
        RECT  0.45 5.15 2.95 5.65 ;
        RECT  1.40 6.65 4.15 7.15 ;
        RECT  3.65 3.85 4.15 8.20 ;
        RECT  3.65 3.85 4.85 4.55 ;
        RECT  4.15 7.70 4.85 9.30 ;
        RECT  4.60 6.25 5.30 7.25 ;
        RECT  4.60 6.75 8.35 7.25 ;
        RECT  7.85 3.95 8.35 9.10 ;
        RECT  7.85 3.95 8.55 4.65 ;
        RECT  7.85 7.50 8.55 9.10 ;
        RECT  8.85 2.45 9.55 3.15 ;
        RECT  8.80 5.45 9.55 6.15 ;
        RECT  9.05 2.45 9.55 10.55 ;
        RECT  8.95 9.85 10.60 10.55 ;
        RECT  10.40 2.75 11.10 4.45 ;
        RECT  10.40 3.95 12.10 4.45 ;
        RECT  11.60 3.95 12.10 8.25 ;
        RECT  11.40 7.55 12.10 8.25 ;
        RECT  11.60 5.65 13.85 6.15 ;
        RECT  13.15 5.65 13.85 6.35 ;
    END
END LGCPX4
MACRO LGCPX8
    CLASS CORE ;
    FOREIGN LGCPX8 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  15.80 2.75 16.50 4.45 ;
        RECT  16.00 2.75 16.50 10.55 ;
        RECT  15.80 7.15 16.50 10.55 ;
        RECT  16.00 5.40 19.35 5.90 ;
        RECT  18.50 2.75 19.00 10.55 ;
        RECT  18.50 2.75 19.20 4.45 ;
        RECT  18.50 7.15 19.20 10.55 ;
        RECT  18.45 5.40 19.35 6.30 ;
        END
    END GCLK
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.85 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END CLK
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.70 2.50 11.00 ;
        RECT  0.45 10.25 2.50 11.00 ;
        RECT  6.50 7.70 7.20 11.00 ;
        RECT  8.30 10.30 10.95 11.00 ;
        RECT  11.75 7.30 12.45 11.00 ;
        RECT  14.45 7.30 15.15 11.00 ;
        RECT  17.15 7.30 17.85 11.00 ;
        RECT  19.85 7.30 20.55 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.50 ;
        RECT  6.50 2.00 7.20 4.65 ;
        RECT  8.90 2.00 9.60 3.05 ;
        RECT  14.30 2.00 15.00 4.45 ;
        RECT  17.15 2.00 17.85 4.45 ;
        RECT  19.85 2.00 20.55 4.45 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.65 7.70 4.85 8.20 ;
        RECT  0.45 3.80 0.95 9.30 ;
        RECT  0.45 3.80 1.15 4.50 ;
        RECT  0.45 7.70 1.15 9.30 ;
        RECT  1.40 6.45 2.10 7.15 ;
        RECT  2.25 4.95 2.95 5.65 ;
        RECT  0.45 5.15 2.95 5.65 ;
        RECT  1.40 6.65 4.15 7.15 ;
        RECT  3.65 3.85 4.15 8.20 ;
        RECT  3.65 3.85 4.85 4.55 ;
        RECT  4.15 7.70 4.85 9.30 ;
        RECT  4.60 6.25 5.30 7.25 ;
        RECT  4.60 6.75 8.35 7.25 ;
        RECT  7.85 3.95 8.35 9.20 ;
        RECT  7.85 3.95 8.55 4.65 ;
        RECT  7.85 7.60 8.55 9.20 ;
        RECT  8.80 5.45 10.75 6.15 ;
        RECT  10.25 2.45 10.75 8.80 ;
        RECT  10.25 2.45 10.95 3.15 ;
        RECT  10.25 7.20 10.95 8.80 ;
        RECT  11.80 2.85 12.50 4.45 ;
        RECT  11.80 3.95 13.80 4.45 ;
        RECT  13.30 3.95 13.80 10.55 ;
        RECT  13.10 7.15 13.80 10.55 ;
        RECT  13.30 5.65 15.55 6.15 ;
        RECT  14.85 5.65 15.55 6.35 ;
    END
END LGCPX8
MACRO LOGIC0
    CLASS CORE ;
    FOREIGN LOGIC0 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  2.05 7.80 2.55 10.20 ;
        RECT  1.65 9.30 2.55 10.20 ;
        RECT  2.95 7.60 3.65 8.30 ;
        RECT  2.05 7.80 3.65 8.30 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.00 11.00 4.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.55 2.00 1.25 8.30 ;
        RECT  0.00 0.00 4.20 2.00 ;
        END
    END gnd!
END LOGIC0
MACRO LOGIC1
    CLASS CORE ;
    FOREIGN LOGIC1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.05 2.85 1.55 7.80 ;
        RECT  0.25 6.65 1.55 7.80 ;
        RECT  1.05 2.85 1.75 3.55 ;
        RECT  0.25 7.10 1.75 7.80 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.05 9.50 1.75 11.00 ;
        RECT  0.00 11.00 2.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.00 0.00 2.80 2.00 ;
        END
    END gnd!
END LOGIC1
MACRO LSGCNX1
    CLASS CORE ;
    FOREIGN LSGCNX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END SE
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.35 1.15 6.35 ;
        RECT  0.45 3.75 1.15 8.70 ;
        END
    END GCLK
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  17.95 5.40 19.35 6.30 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.80 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END CLK
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.95 7.40 2.65 11.00 ;
        RECT  7.35 7.15 7.85 11.00 ;
        RECT  7.35 7.15 8.05 8.75 ;
        RECT  6.35 10.00 8.95 11.00 ;
        RECT  12.45 7.30 13.15 11.00 ;
        RECT  17.15 7.70 18.05 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.40 ;
        RECT  4.50 2.00 5.20 4.40 ;
        RECT  7.35 2.00 8.05 4.40 ;
        RECT  12.45 2.00 13.15 4.05 ;
        RECT  17.15 2.00 17.85 4.00 ;
        RECT  19.85 2.00 20.55 4.00 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.60 6.75 5.05 6.95 ;
        RECT  1.60 4.85 2.10 6.95 ;
        RECT  1.60 6.05 2.30 6.95 ;
        RECT  3.10 6.45 3.60 7.25 ;
        RECT  1.60 6.45 3.60 6.95 ;
        RECT  3.15 3.75 3.85 5.35 ;
        RECT  1.60 4.85 3.85 5.35 ;
        RECT  3.10 6.75 5.05 7.25 ;
        RECT  4.35 6.75 5.05 10.55 ;
        RECT  6.00 3.75 6.70 8.90 ;
        RECT  7.75 6.00 8.45 6.70 ;
        RECT  6.00 6.20 8.45 6.70 ;
        RECT  8.95 3.75 9.45 8.70 ;
        RECT  8.75 7.10 9.45 8.70 ;
        RECT  9.10 2.45 9.80 3.15 ;
        RECT  8.75 3.75 10.60 4.45 ;
        RECT  8.75 8.00 10.60 8.70 ;
        RECT  9.10 2.65 11.60 3.15 ;
        RECT  11.10 2.65 11.60 8.85 ;
        RECT  11.10 3.35 11.80 4.05 ;
        RECT  11.10 7.25 11.80 8.85 ;
        RECT  12.05 6.05 12.75 6.80 ;
        RECT  11.10 4.80 13.55 5.30 ;
        RECT  12.85 4.80 13.55 5.50 ;
        RECT  12.05 6.30 15.50 6.80 ;
        RECT  14.80 3.35 15.50 8.70 ;
        RECT  16.70 5.55 17.40 6.25 ;
        RECT  16.90 4.45 17.40 7.25 ;
        RECT  18.50 3.40 19.00 4.95 ;
        RECT  16.90 4.45 19.00 4.95 ;
        RECT  18.50 3.40 19.20 4.10 ;
        RECT  16.90 6.75 20.40 7.25 ;
        RECT  19.70 6.75 20.40 10.55 ;
    END
END LSGCNX1
MACRO LSGCNX2
    CLASS CORE ;
    FOREIGN LSGCNX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END SE
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.35 1.15 6.35 ;
        RECT  0.45 2.70 1.15 10.55 ;
        END
    END GCLK
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  17.95 5.40 19.35 6.30 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.80 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END CLK
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.90 7.40 2.60 11.00 ;
        RECT  7.35 7.15 7.85 11.00 ;
        RECT  7.35 7.15 8.05 8.75 ;
        RECT  6.35 10.00 8.95 11.00 ;
        RECT  12.45 7.30 13.15 11.00 ;
        RECT  17.15 7.70 18.05 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.40 ;
        RECT  4.65 2.00 5.35 4.40 ;
        RECT  7.50 2.00 8.20 4.40 ;
        RECT  12.45 2.00 13.15 4.05 ;
        RECT  17.15 2.00 17.85 4.00 ;
        RECT  19.85 2.00 20.55 4.00 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.60 6.75 5.05 6.95 ;
        RECT  1.60 4.85 2.10 6.95 ;
        RECT  1.60 6.05 2.30 6.95 ;
        RECT  3.10 6.45 3.60 7.25 ;
        RECT  1.60 6.45 3.60 6.95 ;
        RECT  3.30 3.75 3.80 5.35 ;
        RECT  1.60 4.85 3.80 5.35 ;
        RECT  3.30 3.75 4.00 4.50 ;
        RECT  3.10 6.75 5.05 7.25 ;
        RECT  4.35 6.75 5.05 10.55 ;
        RECT  6.15 3.75 6.70 8.90 ;
        RECT  6.00 7.15 6.70 8.90 ;
        RECT  6.15 3.75 6.85 4.50 ;
        RECT  7.85 6.00 8.55 6.70 ;
        RECT  6.15 6.20 8.55 6.70 ;
        RECT  9.00 3.75 9.50 8.75 ;
        RECT  8.75 7.15 9.50 8.75 ;
        RECT  9.25 2.45 9.95 3.15 ;
        RECT  8.75 8.00 10.60 8.75 ;
        RECT  8.90 3.75 10.65 4.45 ;
        RECT  9.25 2.65 11.60 3.15 ;
        RECT  11.10 2.65 11.60 8.85 ;
        RECT  11.10 3.35 11.80 4.05 ;
        RECT  11.10 7.25 11.80 8.85 ;
        RECT  12.05 6.05 12.75 6.80 ;
        RECT  11.10 4.80 13.55 5.30 ;
        RECT  12.85 4.80 13.55 5.50 ;
        RECT  12.05 6.30 15.50 6.80 ;
        RECT  14.80 3.35 15.50 8.70 ;
        RECT  16.70 5.55 17.40 6.25 ;
        RECT  16.90 4.45 17.40 7.25 ;
        RECT  18.50 3.40 19.00 4.95 ;
        RECT  16.90 4.45 19.00 4.95 ;
        RECT  18.50 3.40 19.20 4.10 ;
        RECT  16.90 6.75 20.40 7.25 ;
        RECT  19.70 6.75 20.40 10.55 ;
    END
END LSGCNX2
MACRO LSGCNX3
    CLASS CORE ;
    FOREIGN LSGCNX3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  21.25 5.40 22.15 6.30 ;
        END
    END SE
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.35 2.55 6.35 ;
        RECT  1.85 3.75 2.55 9.65 ;
        END
    END GCLK
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  19.35 5.40 20.75 6.30 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.80 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END CLK
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 7.40 1.20 11.00 ;
        RECT  0.50 10.90 2.30 11.00 ;
        RECT  3.35 7.40 4.05 11.00 ;
        RECT  8.75 7.15 9.25 11.00 ;
        RECT  8.75 7.15 9.45 8.75 ;
        RECT  7.75 10.00 10.35 11.00 ;
        RECT  13.85 7.30 14.55 11.00 ;
        RECT  18.55 7.70 19.45 11.00 ;
        RECT  0.00 11.00 22.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 2.00 1.20 4.40 ;
        RECT  3.20 2.00 3.90 4.40 ;
        RECT  6.05 2.00 6.75 4.40 ;
        RECT  8.90 2.00 9.60 4.40 ;
        RECT  13.85 2.00 14.55 4.05 ;
        RECT  18.55 2.00 19.25 4.00 ;
        RECT  21.25 2.00 21.95 4.00 ;
        RECT  0.00 0.00 22.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.00 6.75 6.45 6.95 ;
        RECT  3.00 4.85 3.50 6.95 ;
        RECT  3.00 6.05 3.70 6.95 ;
        RECT  4.50 6.45 5.00 7.25 ;
        RECT  3.00 6.45 5.00 6.95 ;
        RECT  4.70 3.75 5.20 5.35 ;
        RECT  3.00 4.85 5.20 5.35 ;
        RECT  4.70 3.75 5.40 4.50 ;
        RECT  4.50 6.75 6.45 7.25 ;
        RECT  5.75 6.75 6.45 10.55 ;
        RECT  7.55 3.75 8.10 8.90 ;
        RECT  7.40 7.15 8.10 8.90 ;
        RECT  7.55 3.75 8.25 4.50 ;
        RECT  9.25 6.00 9.95 6.70 ;
        RECT  7.55 6.20 9.95 6.70 ;
        RECT  10.40 3.75 10.90 8.75 ;
        RECT  10.15 7.15 10.90 8.75 ;
        RECT  10.65 2.45 11.35 3.15 ;
        RECT  10.15 8.00 12.00 8.75 ;
        RECT  10.30 3.75 12.05 4.45 ;
        RECT  10.65 2.65 13.00 3.15 ;
        RECT  12.50 2.65 13.00 8.85 ;
        RECT  12.50 3.35 13.20 4.05 ;
        RECT  12.50 7.25 13.20 8.85 ;
        RECT  13.45 6.05 14.15 6.80 ;
        RECT  12.50 4.80 14.95 5.30 ;
        RECT  14.25 4.80 14.95 5.50 ;
        RECT  13.45 6.30 16.90 6.80 ;
        RECT  16.20 3.35 16.90 8.70 ;
        RECT  18.10 5.55 18.80 6.25 ;
        RECT  18.30 4.45 18.80 7.25 ;
        RECT  19.90 3.40 20.40 4.95 ;
        RECT  18.30 4.45 20.40 4.95 ;
        RECT  19.90 3.40 20.60 4.10 ;
        RECT  18.30 6.75 21.80 7.25 ;
        RECT  21.10 6.75 21.80 10.55 ;
    END
END LSGCNX3
MACRO LSGCNX4
    CLASS CORE ;
    FOREIGN LSGCNX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  21.25 5.40 22.15 6.30 ;
        END
    END SE
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.35 2.55 6.35 ;
        RECT  1.85 2.70 2.55 10.55 ;
        END
    END GCLK
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  19.35 5.40 20.75 6.30 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.80 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END CLK
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 7.40 1.20 11.00 ;
        RECT  3.35 7.40 4.05 11.00 ;
        RECT  8.75 7.15 9.25 11.00 ;
        RECT  8.75 7.15 9.45 8.75 ;
        RECT  7.75 10.00 10.35 11.00 ;
        RECT  13.85 7.30 14.55 11.00 ;
        RECT  18.55 7.70 19.45 11.00 ;
        RECT  0.00 11.00 22.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 2.00 1.20 4.40 ;
        RECT  3.20 2.00 3.90 4.40 ;
        RECT  6.05 2.00 6.75 4.40 ;
        RECT  8.90 2.00 9.60 4.40 ;
        RECT  13.85 2.00 14.55 4.05 ;
        RECT  18.55 2.00 19.25 4.00 ;
        RECT  21.25 2.00 21.95 4.00 ;
        RECT  0.00 0.00 22.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.00 6.75 6.45 6.95 ;
        RECT  3.00 4.85 3.50 6.95 ;
        RECT  3.00 6.05 3.70 6.95 ;
        RECT  4.50 6.45 5.00 7.25 ;
        RECT  3.00 6.45 5.00 6.95 ;
        RECT  4.70 3.75 5.20 5.35 ;
        RECT  3.00 4.85 5.20 5.35 ;
        RECT  4.70 3.75 5.40 4.50 ;
        RECT  4.50 6.75 6.45 7.25 ;
        RECT  5.75 6.75 6.45 10.55 ;
        RECT  7.55 3.75 8.10 8.90 ;
        RECT  7.40 7.15 8.10 8.90 ;
        RECT  7.55 3.75 8.25 4.50 ;
        RECT  9.25 6.00 9.95 6.70 ;
        RECT  7.55 6.20 9.95 6.70 ;
        RECT  10.40 3.75 10.90 8.75 ;
        RECT  10.15 7.15 10.90 8.75 ;
        RECT  10.65 2.45 11.35 3.15 ;
        RECT  10.15 8.00 12.00 8.75 ;
        RECT  10.30 3.75 12.05 4.45 ;
        RECT  10.65 2.65 13.00 3.15 ;
        RECT  12.50 2.65 13.00 8.85 ;
        RECT  12.50 3.35 13.20 4.05 ;
        RECT  12.50 7.25 13.20 8.85 ;
        RECT  13.45 6.05 14.15 6.80 ;
        RECT  12.50 4.80 14.95 5.30 ;
        RECT  14.25 4.80 14.95 5.50 ;
        RECT  13.45 6.30 16.90 6.80 ;
        RECT  16.20 3.35 16.90 8.70 ;
        RECT  18.10 5.55 18.80 6.25 ;
        RECT  18.30 4.45 18.80 7.25 ;
        RECT  19.90 3.40 20.40 4.95 ;
        RECT  18.30 4.45 20.40 4.95 ;
        RECT  19.90 3.40 20.60 4.10 ;
        RECT  18.30 6.75 21.80 7.25 ;
        RECT  21.10 6.75 21.80 10.55 ;
    END
END LSGCNX4
MACRO LSGCNX8
    CLASS CORE ;
    FOREIGN LSGCNX8 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 26.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  25.45 5.40 26.35 6.30 ;
        END
    END SE
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.45 1.15 4.50 ;
        RECT  0.65 2.45 1.15 10.55 ;
        RECT  0.45 7.10 1.15 10.55 ;
        RECT  1.65 5.35 2.55 6.35 ;
        RECT  0.65 5.35 2.55 5.85 ;
        RECT  1.65 5.85 3.65 6.35 ;
        RECT  3.15 2.45 3.65 10.55 ;
        RECT  3.15 2.45 3.85 4.50 ;
        RECT  3.15 7.10 3.85 10.55 ;
        END
    END GCLK
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  23.55 5.40 24.95 6.30 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.55 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END CLK
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.10 2.50 11.00 ;
        RECT  4.50 7.20 5.20 11.00 ;
        RECT  4.50 9.40 8.30 11.00 ;
        RECT  12.95 7.15 13.45 11.00 ;
        RECT  12.95 7.15 13.65 8.75 ;
        RECT  11.95 10.00 14.55 11.00 ;
        RECT  18.05 7.30 18.75 11.00 ;
        RECT  22.75 7.70 23.65 11.00 ;
        RECT  0.00 11.00 26.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.50 ;
        RECT  4.50 2.00 5.20 4.50 ;
        RECT  6.00 2.00 6.70 4.50 ;
        RECT  7.55 2.00 8.25 4.40 ;
        RECT  10.25 2.00 10.95 4.40 ;
        RECT  13.10 2.00 13.80 4.40 ;
        RECT  18.05 2.00 18.75 4.05 ;
        RECT  22.75 2.00 23.45 4.00 ;
        RECT  25.45 2.00 26.15 4.00 ;
        RECT  0.00 0.00 26.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.15 6.05 4.85 6.75 ;
        RECT  4.15 6.25 7.35 6.75 ;
        RECT  6.85 6.25 7.35 7.80 ;
        RECT  8.90 2.70 9.40 7.80 ;
        RECT  8.90 2.70 9.60 4.50 ;
        RECT  6.85 7.10 10.65 7.80 ;
        RECT  9.95 7.10 10.65 10.55 ;
        RECT  11.75 3.75 12.30 8.90 ;
        RECT  11.60 7.15 12.30 8.90 ;
        RECT  11.75 3.75 12.45 4.50 ;
        RECT  13.45 6.00 14.15 6.70 ;
        RECT  11.75 6.20 14.15 6.70 ;
        RECT  14.60 3.75 15.10 8.75 ;
        RECT  14.35 7.15 15.10 8.75 ;
        RECT  14.85 2.45 15.55 3.15 ;
        RECT  14.35 8.00 16.20 8.75 ;
        RECT  14.50 3.75 16.25 4.45 ;
        RECT  14.85 2.65 17.20 3.15 ;
        RECT  16.70 2.65 17.20 8.85 ;
        RECT  16.70 3.35 17.40 4.05 ;
        RECT  16.70 7.25 17.40 8.85 ;
        RECT  17.65 6.05 18.35 6.80 ;
        RECT  16.70 4.80 19.15 5.30 ;
        RECT  18.45 4.80 19.15 5.50 ;
        RECT  17.65 6.30 21.10 6.80 ;
        RECT  20.40 3.35 21.10 8.70 ;
        RECT  22.30 5.55 23.00 6.25 ;
        RECT  22.50 4.45 23.00 7.25 ;
        RECT  24.10 3.40 24.60 4.95 ;
        RECT  22.50 4.45 24.60 4.95 ;
        RECT  24.10 3.40 24.80 4.10 ;
        RECT  22.50 6.75 26.00 7.25 ;
        RECT  25.30 6.75 26.00 10.55 ;
    END
END LSGCNX8
MACRO LSGCPX1
    CLASS CORE ;
    FOREIGN LSGCPX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END SE
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.45 3.35 1.15 4.45 ;
        RECT  0.25 5.35 1.15 6.35 ;
        RECT  0.65 3.35 1.15 8.75 ;
        RECT  0.45 7.10 1.15 8.75 ;
        END
    END GCLK
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.40 19.35 6.30 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END CLK
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.00 ;
        RECT  8.10 2.00 8.80 4.40 ;
        RECT  12.45 2.00 13.15 4.05 ;
        RECT  17.15 2.00 17.85 4.00 ;
        RECT  19.85 2.00 20.55 4.00 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.20 2.50 11.00 ;
        RECT  3.45 9.05 5.35 11.00 ;
        RECT  4.65 7.15 5.35 11.00 ;
        RECT  0.70 10.05 5.35 11.00 ;
        RECT  7.60 7.15 8.10 11.00 ;
        RECT  7.60 7.15 8.30 8.75 ;
        RECT  0.70 10.10 8.85 11.00 ;
        RECT  12.60 7.80 13.30 11.00 ;
        RECT  17.50 8.00 18.20 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    OBS
        LAYER M1M ;
        RECT  9.20 9.25 10.10 9.70 ;
        RECT  1.60 6.05 2.30 6.75 ;
        RECT  1.60 6.20 3.90 6.75 ;
        RECT  3.40 4.45 3.90 7.85 ;
        RECT  3.30 6.20 3.90 7.85 ;
        RECT  3.30 7.15 4.00 7.85 ;
        RECT  4.30 3.40 5.00 4.95 ;
        RECT  3.40 4.45 5.00 4.95 ;
        RECT  6.75 3.75 7.45 4.45 ;
        RECT  6.45 5.95 6.95 8.90 ;
        RECT  6.25 7.15 6.95 8.90 ;
        RECT  6.95 3.75 7.45 6.50 ;
        RECT  6.45 5.95 8.65 6.50 ;
        RECT  7.95 5.95 8.65 6.70 ;
        RECT  8.95 7.15 9.70 8.75 ;
        RECT  9.45 3.80 9.70 9.95 ;
        RECT  9.20 5.85 9.70 9.70 ;
        RECT  9.45 3.80 9.95 6.30 ;
        RECT  9.20 5.85 9.95 6.30 ;
        RECT  9.40 9.25 10.10 9.95 ;
        RECT  9.45 3.80 10.20 4.50 ;
        RECT  11.10 3.40 11.60 9.35 ;
        RECT  11.10 3.40 11.80 4.10 ;
        RECT  11.10 7.75 11.95 9.35 ;
        RECT  11.10 5.30 13.55 5.80 ;
        RECT  12.20 6.55 12.90 7.30 ;
        RECT  12.85 5.30 13.55 6.00 ;
        RECT  12.20 6.80 15.65 7.30 ;
        RECT  14.45 3.35 14.95 7.30 ;
        RECT  14.50 9.75 15.20 10.45 ;
        RECT  14.45 3.35 15.50 4.05 ;
        RECT  14.95 6.80 15.65 9.20 ;
        RECT  15.40 4.70 16.60 5.40 ;
        RECT  16.10 4.70 16.60 10.45 ;
        RECT  14.50 9.95 16.60 10.45 ;
        RECT  17.15 4.45 17.65 7.25 ;
        RECT  17.15 5.50 17.85 6.20 ;
        RECT  18.50 3.40 19.00 4.95 ;
        RECT  17.15 4.45 19.00 4.95 ;
        RECT  18.50 3.40 19.20 4.10 ;
        RECT  17.15 6.75 20.55 7.25 ;
        RECT  19.85 6.75 20.55 10.55 ;
    END
END LSGCPX1
MACRO LSGCPX2
    CLASS CORE ;
    FOREIGN LSGCPX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END SE
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.50 1.15 4.45 ;
        RECT  0.25 5.35 1.15 6.35 ;
        RECT  0.65 2.50 1.15 10.55 ;
        RECT  0.45 7.10 1.15 10.55 ;
        END
    END GCLK
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.40 19.35 6.30 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END CLK
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 3.90 ;
        RECT  8.10 2.00 8.80 4.40 ;
        RECT  12.45 2.00 13.15 4.05 ;
        RECT  17.15 2.00 17.85 4.00 ;
        RECT  19.85 2.00 20.55 4.00 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.25 2.50 11.00 ;
        RECT  4.65 7.15 5.35 11.00 ;
        RECT  3.45 9.05 5.35 11.00 ;
        RECT  7.60 7.15 8.10 11.00 ;
        RECT  7.60 7.15 8.30 8.75 ;
        RECT  3.45 10.10 8.85 11.00 ;
        RECT  12.60 7.80 13.30 11.00 ;
        RECT  17.50 8.00 18.20 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    OBS
        LAYER M1M ;
        RECT  9.20 9.25 10.10 9.70 ;
        RECT  1.60 6.05 2.30 6.75 ;
        RECT  1.60 6.20 3.90 6.75 ;
        RECT  3.40 4.45 3.90 7.85 ;
        RECT  3.30 6.20 3.90 7.85 ;
        RECT  3.30 7.15 4.00 7.85 ;
        RECT  4.30 3.40 5.00 4.95 ;
        RECT  3.40 4.45 5.00 4.95 ;
        RECT  6.75 3.75 7.45 4.45 ;
        RECT  6.45 5.95 6.95 8.90 ;
        RECT  6.25 7.15 6.95 8.90 ;
        RECT  6.95 3.75 7.45 6.50 ;
        RECT  6.45 5.95 8.65 6.50 ;
        RECT  7.95 5.95 8.65 6.70 ;
        RECT  8.95 7.15 9.70 8.75 ;
        RECT  9.45 3.80 9.70 9.95 ;
        RECT  9.20 5.85 9.70 9.70 ;
        RECT  9.45 3.80 9.95 6.30 ;
        RECT  9.20 5.85 9.95 6.30 ;
        RECT  9.40 9.25 10.10 9.95 ;
        RECT  9.45 3.80 10.20 4.50 ;
        RECT  11.10 3.40 11.60 9.35 ;
        RECT  11.10 3.40 11.80 4.10 ;
        RECT  11.10 7.75 11.95 9.35 ;
        RECT  11.10 5.30 13.55 5.80 ;
        RECT  12.20 6.55 12.90 7.30 ;
        RECT  12.85 5.30 13.55 6.00 ;
        RECT  12.20 6.80 15.65 7.30 ;
        RECT  14.45 3.35 14.95 7.30 ;
        RECT  14.50 9.75 15.20 10.45 ;
        RECT  14.45 3.35 15.50 4.05 ;
        RECT  14.95 6.80 15.65 9.20 ;
        RECT  15.40 4.70 16.60 5.40 ;
        RECT  16.10 4.70 16.60 10.45 ;
        RECT  14.50 9.95 16.60 10.45 ;
        RECT  17.15 4.45 17.65 7.25 ;
        RECT  17.15 5.50 17.85 6.20 ;
        RECT  18.50 3.40 19.00 4.95 ;
        RECT  17.15 4.45 19.00 4.95 ;
        RECT  18.50 3.40 19.20 4.10 ;
        RECT  17.15 6.75 20.55 7.25 ;
        RECT  19.85 6.75 20.55 10.55 ;
    END
END LSGCPX2
MACRO LSGCPX3
    CLASS CORE ;
    FOREIGN LSGCPX3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  21.25 5.40 22.15 6.30 ;
        END
    END SE
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.35 1.15 6.35 ;
        RECT  0.25 5.65 2.45 6.15 ;
        RECT  1.95 4.45 2.45 9.40 ;
        RECT  1.95 7.10 2.65 9.40 ;
        RECT  2.50 3.15 3.00 4.95 ;
        RECT  1.95 4.45 3.00 4.95 ;
        RECT  2.50 3.15 3.20 3.85 ;
        END
    END GCLK
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END CLK
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.15 2.00 1.85 3.85 ;
        RECT  4.00 2.00 4.70 4.00 ;
        RECT  9.50 2.00 10.20 4.40 ;
        RECT  13.85 2.00 14.55 4.05 ;
        RECT  18.55 2.00 19.25 4.00 ;
        RECT  21.25 2.00 21.95 4.00 ;
        RECT  0.00 0.00 22.40 2.00 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.60 7.10 1.30 11.00 ;
        RECT  3.30 7.25 4.00 11.00 ;
        RECT  6.15 7.15 6.85 11.00 ;
        RECT  9.00 7.15 9.50 11.00 ;
        RECT  9.00 7.15 9.70 8.75 ;
        RECT  4.85 10.10 10.25 11.00 ;
        RECT  14.00 7.80 14.70 11.00 ;
        RECT  18.90 8.00 19.60 11.00 ;
        RECT  0.00 11.00 22.40 13.00 ;
        END
    END vdd!
    OBS
        LAYER M1M ;
        RECT  10.60 9.25 11.50 9.70 ;
        RECT  3.10 6.05 3.80 6.75 ;
        RECT  3.10 6.20 5.30 6.75 ;
        RECT  4.80 4.45 5.30 8.75 ;
        RECT  4.80 7.15 5.50 8.75 ;
        RECT  6.35 2.55 7.05 4.95 ;
        RECT  4.80 4.45 7.05 4.95 ;
        RECT  8.15 3.75 8.85 4.45 ;
        RECT  7.85 5.95 8.35 8.90 ;
        RECT  7.65 7.15 8.35 8.90 ;
        RECT  8.35 3.75 8.85 6.50 ;
        RECT  7.85 5.95 10.05 6.50 ;
        RECT  9.35 5.95 10.05 6.70 ;
        RECT  10.35 7.15 11.10 8.75 ;
        RECT  10.85 3.80 11.10 9.95 ;
        RECT  10.60 5.85 11.10 9.70 ;
        RECT  10.85 3.80 11.35 6.30 ;
        RECT  10.60 5.85 11.35 6.30 ;
        RECT  10.80 9.25 11.50 9.95 ;
        RECT  10.85 3.80 11.60 4.50 ;
        RECT  12.50 3.40 13.00 9.35 ;
        RECT  12.50 3.40 13.20 4.10 ;
        RECT  12.50 7.75 13.35 9.35 ;
        RECT  12.50 5.30 14.95 5.80 ;
        RECT  13.60 6.55 14.30 7.30 ;
        RECT  14.25 5.30 14.95 6.00 ;
        RECT  13.60 6.80 17.05 7.30 ;
        RECT  15.85 3.35 16.35 7.30 ;
        RECT  15.90 9.75 16.60 10.45 ;
        RECT  15.85 3.35 16.90 4.05 ;
        RECT  16.35 6.80 17.05 9.20 ;
        RECT  16.80 4.70 18.00 5.40 ;
        RECT  17.50 4.70 18.00 10.45 ;
        RECT  15.90 9.95 18.00 10.45 ;
        RECT  18.55 4.45 19.05 7.25 ;
        RECT  18.55 5.50 19.25 6.20 ;
        RECT  19.90 3.40 20.40 4.95 ;
        RECT  18.55 4.45 20.40 4.95 ;
        RECT  19.90 3.40 20.60 4.10 ;
        RECT  18.55 6.75 21.95 7.25 ;
        RECT  21.25 6.75 21.95 10.55 ;
    END
END LSGCPX3
MACRO LSGCPX4
    CLASS CORE ;
    FOREIGN LSGCPX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  21.25 5.40 22.15 6.30 ;
        END
    END SE
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.35 1.15 6.35 ;
        RECT  0.25 5.65 2.45 6.15 ;
        RECT  1.95 4.45 2.45 10.55 ;
        RECT  1.95 7.10 2.65 10.55 ;
        RECT  2.65 2.55 3.15 4.95 ;
        RECT  1.95 4.45 3.15 4.95 ;
        RECT  2.65 2.55 3.35 4.55 ;
        RECT  1.95 4.45 3.35 4.55 ;
        END
    END GCLK
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END CLK
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.30 2.00 2.00 4.00 ;
        RECT  4.00 2.00 4.70 4.00 ;
        RECT  9.50 2.00 10.20 4.40 ;
        RECT  13.85 2.00 14.55 4.05 ;
        RECT  18.55 2.00 19.25 4.00 ;
        RECT  21.25 2.00 21.95 4.00 ;
        RECT  0.00 0.00 22.40 2.00 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.60 7.10 1.30 11.00 ;
        RECT  3.30 7.25 4.00 11.00 ;
        RECT  6.15 7.15 6.85 11.00 ;
        RECT  9.00 7.15 9.50 11.00 ;
        RECT  9.00 7.15 9.70 8.75 ;
        RECT  4.85 10.10 10.25 11.00 ;
        RECT  14.00 7.80 14.70 11.00 ;
        RECT  18.90 8.00 19.60 11.00 ;
        RECT  0.00 11.00 22.40 13.00 ;
        END
    END vdd!
    OBS
        LAYER M1M ;
        RECT  10.60 9.25 11.50 9.70 ;
        RECT  3.10 6.05 3.80 6.75 ;
        RECT  3.10 6.20 5.30 6.75 ;
        RECT  4.80 4.45 5.30 8.75 ;
        RECT  4.80 7.15 5.50 8.75 ;
        RECT  6.35 2.55 7.05 4.95 ;
        RECT  4.80 4.45 7.05 4.95 ;
        RECT  8.15 3.75 8.85 4.45 ;
        RECT  7.85 5.95 8.35 8.90 ;
        RECT  7.65 7.15 8.35 8.90 ;
        RECT  8.35 3.75 8.85 6.50 ;
        RECT  7.85 5.95 10.05 6.50 ;
        RECT  9.35 5.95 10.05 6.70 ;
        RECT  10.35 7.15 11.10 8.75 ;
        RECT  10.85 3.80 11.10 9.95 ;
        RECT  10.60 5.85 11.10 9.70 ;
        RECT  10.85 3.80 11.35 6.30 ;
        RECT  10.60 5.85 11.35 6.30 ;
        RECT  10.80 9.25 11.50 9.95 ;
        RECT  10.85 3.80 11.60 4.50 ;
        RECT  12.50 3.40 13.00 9.35 ;
        RECT  12.50 3.40 13.20 4.10 ;
        RECT  12.50 7.75 13.35 9.35 ;
        RECT  12.50 5.30 14.95 5.80 ;
        RECT  13.60 6.55 14.30 7.30 ;
        RECT  14.25 5.30 14.95 6.00 ;
        RECT  13.60 6.80 17.05 7.30 ;
        RECT  15.85 3.35 16.35 7.30 ;
        RECT  15.90 9.75 16.60 10.45 ;
        RECT  15.85 3.35 16.90 4.05 ;
        RECT  16.35 6.80 17.05 9.20 ;
        RECT  16.80 4.70 18.00 5.40 ;
        RECT  17.50 4.70 18.00 10.45 ;
        RECT  15.90 9.95 18.00 10.45 ;
        RECT  18.55 4.45 19.05 7.25 ;
        RECT  18.55 5.50 19.25 6.20 ;
        RECT  19.90 3.40 20.40 4.95 ;
        RECT  18.55 4.45 20.40 4.95 ;
        RECT  19.90 3.40 20.60 4.10 ;
        RECT  18.55 6.75 21.95 7.25 ;
        RECT  21.25 6.75 21.95 10.55 ;
    END
END LSGCPX4
MACRO LSGCPX8
    CLASS CORE ;
    FOREIGN LSGCPX8 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  22.65 5.40 23.55 6.30 ;
        END
    END SE
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.50 1.20 4.55 ;
        RECT  1.00 2.50 1.20 10.55 ;
        RECT  0.70 2.50 1.20 6.10 ;
        RECT  1.00 5.60 1.50 10.55 ;
        RECT  0.80 7.10 1.50 10.55 ;
        RECT  1.65 5.35 2.55 6.35 ;
        RECT  1.00 5.60 2.55 6.35 ;
        RECT  3.15 2.50 3.70 6.60 ;
        RECT  3.15 6.10 4.00 6.60 ;
        RECT  3.50 2.50 3.70 10.55 ;
        RECT  0.70 5.60 3.70 6.10 ;
        RECT  3.15 2.50 3.85 4.50 ;
        RECT  3.50 6.10 4.00 10.55 ;
        RECT  3.50 7.10 4.20 10.55 ;
        END
    END GCLK
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  21.25 5.40 22.15 6.30 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.85 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END CLK
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.50 ;
        RECT  4.50 2.00 5.20 4.50 ;
        RECT  10.90 2.00 11.60 4.40 ;
        RECT  15.25 2.00 15.95 4.05 ;
        RECT  19.95 2.00 20.65 4.00 ;
        RECT  22.65 2.00 23.35 4.00 ;
        RECT  0.00 0.00 23.80 2.00 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.15 7.10 2.85 11.00 ;
        RECT  4.85 7.25 5.55 11.00 ;
        RECT  7.55 7.35 8.25 11.00 ;
        RECT  10.40 7.15 10.90 11.00 ;
        RECT  10.40 7.15 11.10 8.75 ;
        RECT  9.05 10.10 11.65 11.00 ;
        RECT  15.40 7.80 16.10 11.00 ;
        RECT  20.30 8.00 21.00 11.00 ;
        RECT  0.00 11.00 23.80 13.00 ;
        END
    END vdd!
    OBS
        LAYER M1M ;
        RECT  12.00 9.25 12.90 9.70 ;
        RECT  4.15 4.95 4.85 5.65 ;
        RECT  4.15 5.10 6.70 5.65 ;
        RECT  6.20 3.80 6.70 10.55 ;
        RECT  6.20 8.05 6.90 10.55 ;
        RECT  8.00 2.50 8.75 4.50 ;
        RECT  6.20 3.80 8.75 4.50 ;
        RECT  9.55 3.75 10.25 4.45 ;
        RECT  9.25 5.95 9.75 8.90 ;
        RECT  9.05 7.15 9.75 8.90 ;
        RECT  9.75 3.75 10.25 6.50 ;
        RECT  9.25 5.95 11.45 6.50 ;
        RECT  10.75 5.95 11.45 6.70 ;
        RECT  11.75 7.15 12.50 8.75 ;
        RECT  12.25 3.80 12.50 9.95 ;
        RECT  12.00 5.85 12.50 9.70 ;
        RECT  12.25 3.80 12.75 6.30 ;
        RECT  12.00 5.85 12.75 6.30 ;
        RECT  12.20 9.25 12.90 9.95 ;
        RECT  12.25 3.80 13.00 4.50 ;
        RECT  13.90 3.40 14.40 9.35 ;
        RECT  13.90 3.40 14.60 4.10 ;
        RECT  13.90 7.75 14.75 9.35 ;
        RECT  13.90 5.30 16.35 5.80 ;
        RECT  15.00 6.55 15.70 7.30 ;
        RECT  15.65 5.30 16.35 6.00 ;
        RECT  15.00 6.80 18.45 7.30 ;
        RECT  17.25 3.35 17.75 7.30 ;
        RECT  17.30 9.75 18.00 10.45 ;
        RECT  17.25 3.35 18.30 4.05 ;
        RECT  17.75 6.80 18.45 9.20 ;
        RECT  18.20 4.70 19.40 5.40 ;
        RECT  18.90 4.70 19.40 10.45 ;
        RECT  17.30 9.95 19.40 10.45 ;
        RECT  19.95 4.45 20.45 7.25 ;
        RECT  19.95 5.50 20.65 6.20 ;
        RECT  21.30 3.40 21.80 4.95 ;
        RECT  19.95 4.45 21.80 4.95 ;
        RECT  21.30 3.40 22.00 4.10 ;
        RECT  19.95 6.75 23.35 7.25 ;
        RECT  22.65 6.75 23.35 10.55 ;
    END
END LSGCPX8
MACRO LSOGCNX1
    CLASS CORE ;
    FOREIGN LSOGCNX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  21.25 5.40 22.15 6.30 ;
        END
    END SE
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.35 1.15 6.35 ;
        RECT  0.45 3.75 1.15 8.80 ;
        END
    END GCLK
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  19.25 5.40 20.75 6.30 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.80 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END CLK
    PIN CGOBS
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M2M ;
        RECT  12.90 2.70 13.50 8.45 ;
        RECT  12.90 2.70 13.70 3.80 ;
        RECT  12.90 7.35 13.70 8.45 ;
        LAYER M1M ;
        RECT  12.85 2.80 13.80 4.10 ;
        RECT  12.85 7.35 13.80 8.95 ;
        END
    END CGOBS
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 10.05 1.15 11.00 ;
        RECT  1.95 7.40 2.65 11.00 ;
        RECT  7.35 7.15 7.85 11.00 ;
        RECT  7.35 7.15 8.05 8.75 ;
        RECT  6.35 10.00 8.55 11.00 ;
        RECT  11.70 7.35 12.25 11.00 ;
        RECT  11.70 7.35 12.40 8.95 ;
        RECT  14.70 7.30 15.40 11.00 ;
        RECT  19.40 7.75 20.30 11.00 ;
        RECT  0.00 11.00 23.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.40 ;
        RECT  4.65 2.00 5.35 4.40 ;
        RECT  7.50 2.00 8.20 4.40 ;
        RECT  11.70 2.00 12.40 4.05 ;
        RECT  14.70 2.00 15.40 4.10 ;
        RECT  19.40 2.00 20.10 4.00 ;
        RECT  22.10 2.00 22.80 4.00 ;
        RECT  0.00 0.00 23.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.60 6.75 5.05 6.95 ;
        RECT  1.60 4.85 2.10 6.95 ;
        RECT  1.60 6.05 2.30 6.95 ;
        RECT  3.10 6.45 3.60 7.25 ;
        RECT  1.60 6.45 3.60 6.95 ;
        RECT  3.30 3.75 3.80 5.35 ;
        RECT  1.60 4.85 3.80 5.35 ;
        RECT  3.30 3.75 4.00 4.50 ;
        RECT  3.10 6.75 5.05 7.25 ;
        RECT  4.35 6.75 5.05 10.55 ;
        RECT  6.15 3.75 6.70 8.90 ;
        RECT  6.00 7.15 6.70 8.90 ;
        RECT  6.15 3.75 6.85 4.50 ;
        RECT  7.85 6.00 8.55 6.70 ;
        RECT  6.15 6.20 8.55 6.70 ;
        RECT  8.75 7.15 9.50 8.75 ;
        RECT  9.00 3.70 9.50 9.95 ;
        RECT  8.85 3.70 9.55 4.45 ;
        RECT  9.00 9.45 10.70 9.95 ;
        RECT  10.00 9.45 10.70 10.15 ;
        RECT  10.35 3.40 10.85 8.90 ;
        RECT  10.35 7.30 11.05 8.90 ;
        RECT  10.35 3.40 11.10 4.10 ;
        RECT  12.20 6.10 12.90 6.85 ;
        RECT  10.35 5.15 15.80 5.65 ;
        RECT  15.10 5.15 15.80 5.85 ;
        RECT  16.45 3.30 16.95 6.85 ;
        RECT  12.20 6.35 17.55 6.85 ;
        RECT  16.60 9.50 17.30 10.20 ;
        RECT  17.05 6.35 17.55 8.75 ;
        RECT  16.45 3.30 17.75 4.00 ;
        RECT  17.05 7.15 17.75 8.75 ;
        RECT  17.70 4.55 18.70 5.25 ;
        RECT  18.20 4.55 18.70 10.00 ;
        RECT  16.60 9.50 18.70 10.00 ;
        RECT  20.75 3.35 21.45 4.05 ;
        RECT  20.95 3.35 21.45 4.95 ;
        RECT  21.95 7.15 22.65 10.55 ;
        RECT  20.95 4.45 23.25 4.95 ;
        RECT  22.75 4.45 23.25 7.65 ;
        RECT  21.95 7.15 23.25 7.65 ;
        RECT  22.75 5.45 23.45 6.15 ;
        LAYER V1M ;
        RECT  12.80 6.65 13.80 7.65 ;
        RECT  12.80 7.95 13.80 8.95 ;
        RECT  12.80 2.75 13.80 3.75 ;
    END
END LSOGCNX1
MACRO LSOGCNX2
    CLASS CORE ;
    FOREIGN LSOGCNX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  21.25 5.40 22.15 6.30 ;
        END
    END SE
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.35 1.15 6.35 ;
        RECT  0.45 3.40 1.15 10.55 ;
        END
    END GCLK
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  19.25 5.40 20.75 6.30 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.80 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END CLK
    PIN CGOBS
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M2M ;
        RECT  12.90 2.70 13.50 8.45 ;
        RECT  12.90 2.70 13.70 3.80 ;
        RECT  12.90 7.35 13.70 8.45 ;
        LAYER M1M ;
        RECT  12.85 2.80 13.80 4.10 ;
        RECT  12.85 7.35 13.80 8.95 ;
        END
    END CGOBS
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.95 7.40 2.65 11.00 ;
        RECT  7.35 7.15 7.85 11.00 ;
        RECT  7.35 7.15 8.05 8.75 ;
        RECT  6.35 10.00 8.55 11.00 ;
        RECT  11.70 7.35 12.25 11.00 ;
        RECT  11.70 7.35 12.40 8.95 ;
        RECT  14.70 7.30 15.40 11.00 ;
        RECT  19.40 7.75 20.30 11.00 ;
        RECT  0.00 11.00 23.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.05 ;
        RECT  4.65 2.00 5.35 4.40 ;
        RECT  7.50 2.00 8.20 4.40 ;
        RECT  11.70 2.00 12.40 4.05 ;
        RECT  14.70 2.00 15.40 4.10 ;
        RECT  19.40 2.00 20.10 4.00 ;
        RECT  22.10 2.00 22.80 4.00 ;
        RECT  0.00 0.00 23.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.60 6.75 5.05 6.95 ;
        RECT  1.60 4.85 2.10 6.95 ;
        RECT  1.60 6.05 2.30 6.95 ;
        RECT  3.10 6.45 3.60 7.25 ;
        RECT  1.60 6.45 3.60 6.95 ;
        RECT  3.30 3.75 3.80 5.35 ;
        RECT  1.60 4.85 3.80 5.35 ;
        RECT  3.30 3.75 4.00 4.50 ;
        RECT  3.10 6.75 5.05 7.25 ;
        RECT  4.35 6.75 5.05 10.55 ;
        RECT  6.15 3.75 6.70 8.90 ;
        RECT  6.00 7.15 6.70 8.90 ;
        RECT  6.15 3.75 6.85 4.50 ;
        RECT  7.85 6.00 8.55 6.70 ;
        RECT  6.15 6.20 8.55 6.70 ;
        RECT  8.75 7.15 9.50 8.75 ;
        RECT  9.00 3.70 9.50 9.95 ;
        RECT  8.85 3.70 9.55 4.45 ;
        RECT  9.00 9.45 10.70 9.95 ;
        RECT  10.00 9.45 10.70 10.15 ;
        RECT  10.35 3.40 10.85 8.90 ;
        RECT  10.35 7.30 11.05 8.90 ;
        RECT  10.35 3.40 11.10 4.10 ;
        RECT  12.20 6.10 12.90 6.85 ;
        RECT  10.35 5.15 15.80 5.65 ;
        RECT  15.10 5.15 15.80 5.85 ;
        RECT  16.45 3.30 16.95 6.85 ;
        RECT  12.20 6.35 17.55 6.85 ;
        RECT  16.60 9.50 17.30 10.20 ;
        RECT  17.05 6.35 17.55 8.75 ;
        RECT  16.45 3.30 17.75 4.00 ;
        RECT  17.05 7.15 17.75 8.75 ;
        RECT  17.70 4.55 18.70 5.25 ;
        RECT  18.20 4.55 18.70 10.00 ;
        RECT  16.60 9.50 18.70 10.00 ;
        RECT  20.75 3.35 21.45 4.05 ;
        RECT  20.95 3.35 21.45 4.95 ;
        RECT  21.95 7.15 22.65 10.55 ;
        RECT  20.95 4.45 23.25 4.95 ;
        RECT  22.75 4.45 23.25 7.65 ;
        RECT  21.95 7.15 23.25 7.65 ;
        RECT  22.75 5.45 23.45 6.15 ;
        LAYER V1M ;
        RECT  12.80 6.65 13.80 7.65 ;
        RECT  12.80 7.95 13.80 8.95 ;
        RECT  12.80 2.75 13.80 3.75 ;
    END
END LSOGCNX2
MACRO LSOGCNX3
    CLASS CORE ;
    FOREIGN LSOGCNX3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 25.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  22.65 5.40 23.55 6.30 ;
        END
    END SE
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.35 2.55 6.35 ;
        RECT  1.85 3.40 2.55 9.75 ;
        END
    END GCLK
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  20.65 5.40 22.15 6.30 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.80 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END CLK
    PIN CGOBS
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M2M ;
        RECT  14.30 2.70 14.90 8.45 ;
        RECT  14.30 2.70 15.10 3.80 ;
        RECT  14.30 7.35 15.10 8.45 ;
        LAYER M1M ;
        RECT  14.25 2.80 15.20 4.10 ;
        RECT  14.25 7.35 15.20 8.95 ;
        END
    END CGOBS
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 7.40 1.20 11.00 ;
        RECT  3.35 7.40 4.05 11.00 ;
        RECT  8.75 7.15 9.25 11.00 ;
        RECT  8.75 7.15 9.45 8.75 ;
        RECT  7.75 10.00 9.95 11.00 ;
        RECT  13.10 7.35 13.65 11.00 ;
        RECT  13.10 7.35 13.80 8.95 ;
        RECT  16.10 7.30 16.80 11.00 ;
        RECT  20.80 7.75 21.70 11.00 ;
        RECT  0.00 11.00 25.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 2.00 1.20 4.10 ;
        RECT  3.20 2.00 3.90 4.05 ;
        RECT  6.05 2.00 6.75 4.40 ;
        RECT  8.90 2.00 9.60 4.40 ;
        RECT  13.10 2.00 13.80 4.05 ;
        RECT  16.10 2.00 16.80 4.10 ;
        RECT  20.80 2.00 21.50 4.00 ;
        RECT  23.50 2.00 24.20 4.00 ;
        RECT  0.00 0.00 25.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.00 6.75 6.45 6.95 ;
        RECT  3.00 4.85 3.50 6.95 ;
        RECT  3.00 6.05 3.70 6.95 ;
        RECT  4.50 6.45 5.00 7.25 ;
        RECT  3.00 6.45 5.00 6.95 ;
        RECT  4.70 3.75 5.20 5.35 ;
        RECT  3.00 4.85 5.20 5.35 ;
        RECT  4.70 3.75 5.40 4.50 ;
        RECT  4.50 6.75 6.45 7.25 ;
        RECT  5.75 6.75 6.45 10.55 ;
        RECT  7.55 3.75 8.10 8.90 ;
        RECT  7.40 7.15 8.10 8.90 ;
        RECT  7.55 3.75 8.25 4.50 ;
        RECT  9.25 6.00 9.95 6.70 ;
        RECT  7.55 6.20 9.95 6.70 ;
        RECT  10.15 7.15 10.90 8.75 ;
        RECT  10.40 3.70 10.90 9.95 ;
        RECT  10.25 3.70 10.95 4.45 ;
        RECT  10.40 9.45 12.10 9.95 ;
        RECT  11.40 9.45 12.10 10.15 ;
        RECT  11.75 3.40 12.25 8.90 ;
        RECT  11.75 7.30 12.45 8.90 ;
        RECT  11.75 3.40 12.50 4.10 ;
        RECT  13.60 6.10 14.30 6.85 ;
        RECT  11.75 5.15 17.20 5.65 ;
        RECT  16.50 5.15 17.20 5.85 ;
        RECT  17.85 3.30 18.35 6.85 ;
        RECT  13.60 6.35 18.95 6.85 ;
        RECT  18.00 9.50 18.70 10.20 ;
        RECT  18.45 6.35 18.95 8.75 ;
        RECT  17.85 3.30 19.15 4.00 ;
        RECT  18.45 7.15 19.15 8.75 ;
        RECT  19.10 4.55 20.10 5.25 ;
        RECT  19.60 4.55 20.10 10.00 ;
        RECT  18.00 9.50 20.10 10.00 ;
        RECT  22.15 3.35 22.85 4.05 ;
        RECT  22.35 3.35 22.85 4.95 ;
        RECT  23.35 7.15 24.05 10.55 ;
        RECT  22.35 4.45 24.65 4.95 ;
        RECT  24.15 4.45 24.65 7.65 ;
        RECT  23.35 7.15 24.65 7.65 ;
        RECT  24.15 5.45 24.85 6.15 ;
        LAYER V1M ;
        RECT  14.20 6.65 15.20 7.65 ;
        RECT  14.20 7.95 15.20 8.95 ;
        RECT  14.20 2.75 15.20 3.75 ;
    END
END LSOGCNX3
MACRO LSOGCNX4
    CLASS CORE ;
    FOREIGN LSOGCNX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 25.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  22.65 5.40 23.55 6.30 ;
        END
    END SE
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.35 2.55 6.35 ;
        RECT  1.85 2.70 2.55 10.55 ;
        END
    END GCLK
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  20.65 5.40 22.15 6.30 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.80 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END CLK
    PIN CGOBS
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M2M ;
        RECT  14.30 2.70 14.90 8.45 ;
        RECT  14.30 2.70 15.10 3.80 ;
        RECT  14.30 7.35 15.10 8.45 ;
        LAYER M1M ;
        RECT  14.25 2.80 15.20 4.10 ;
        RECT  14.25 7.35 15.20 8.95 ;
        END
    END CGOBS
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 7.40 1.20 11.00 ;
        RECT  3.35 7.40 4.05 11.00 ;
        RECT  8.75 7.15 9.25 11.00 ;
        RECT  8.75 7.15 9.45 8.75 ;
        RECT  7.75 10.00 9.95 11.00 ;
        RECT  13.10 7.35 13.65 11.00 ;
        RECT  13.10 7.35 13.80 8.95 ;
        RECT  16.10 7.30 16.80 11.00 ;
        RECT  20.80 7.75 21.70 11.00 ;
        RECT  0.00 11.00 25.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 2.00 1.20 4.40 ;
        RECT  3.20 2.00 3.90 4.40 ;
        RECT  6.05 2.00 6.75 4.40 ;
        RECT  8.90 2.00 9.60 4.40 ;
        RECT  13.10 2.00 13.80 4.05 ;
        RECT  16.10 2.00 16.80 4.10 ;
        RECT  20.80 2.00 21.50 4.00 ;
        RECT  23.50 2.00 24.20 4.00 ;
        RECT  0.00 0.00 25.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.00 6.75 6.45 6.95 ;
        RECT  3.00 4.85 3.50 6.95 ;
        RECT  3.00 6.05 3.70 6.95 ;
        RECT  4.50 6.45 5.00 7.25 ;
        RECT  3.00 6.45 5.00 6.95 ;
        RECT  4.70 3.75 5.20 5.35 ;
        RECT  3.00 4.85 5.20 5.35 ;
        RECT  4.70 3.75 5.40 4.50 ;
        RECT  4.50 6.75 6.45 7.25 ;
        RECT  5.75 6.75 6.45 10.55 ;
        RECT  7.55 3.75 8.10 8.90 ;
        RECT  7.40 7.15 8.10 8.90 ;
        RECT  7.55 3.75 8.25 4.50 ;
        RECT  9.25 6.00 9.95 6.70 ;
        RECT  7.55 6.20 9.95 6.70 ;
        RECT  10.15 7.15 10.90 8.75 ;
        RECT  10.40 3.70 10.90 9.95 ;
        RECT  10.25 3.70 10.95 4.45 ;
        RECT  10.40 9.45 12.10 9.95 ;
        RECT  11.40 9.45 12.10 10.15 ;
        RECT  11.75 3.40 12.25 8.90 ;
        RECT  11.75 7.30 12.45 8.90 ;
        RECT  11.75 3.40 12.50 4.10 ;
        RECT  13.60 6.10 14.30 6.85 ;
        RECT  11.75 5.15 17.20 5.65 ;
        RECT  16.50 5.15 17.20 5.85 ;
        RECT  17.85 3.30 18.35 6.85 ;
        RECT  13.60 6.35 18.95 6.85 ;
        RECT  18.00 9.50 18.70 10.20 ;
        RECT  18.45 6.35 18.95 8.75 ;
        RECT  17.85 3.30 19.15 4.00 ;
        RECT  18.45 7.15 19.15 8.75 ;
        RECT  19.10 4.55 20.10 5.25 ;
        RECT  19.60 4.55 20.10 10.00 ;
        RECT  18.00 9.50 20.10 10.00 ;
        RECT  22.15 3.35 22.85 4.05 ;
        RECT  22.35 3.35 22.85 4.95 ;
        RECT  23.35 7.15 24.05 10.55 ;
        RECT  22.35 4.45 24.65 4.95 ;
        RECT  24.15 4.45 24.65 7.65 ;
        RECT  23.35 7.15 24.65 7.65 ;
        RECT  24.15 5.45 24.85 6.15 ;
        LAYER V1M ;
        RECT  14.20 6.65 15.20 7.65 ;
        RECT  14.20 7.95 15.20 8.95 ;
        RECT  14.20 2.75 15.20 3.75 ;
    END
END LSOGCNX4
MACRO LSOGCNX8
    CLASS CORE ;
    FOREIGN LSOGCNX8 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 29.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  26.85 5.40 27.75 6.30 ;
        END
    END SE
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.45 1.15 4.50 ;
        RECT  0.65 2.45 1.15 10.55 ;
        RECT  0.45 7.10 1.15 10.55 ;
        RECT  1.65 5.35 2.55 6.35 ;
        RECT  0.65 5.35 2.55 5.85 ;
        RECT  1.65 5.85 3.65 6.35 ;
        RECT  3.15 2.45 3.65 10.55 ;
        RECT  3.15 2.45 3.85 4.50 ;
        RECT  3.15 7.10 3.85 10.55 ;
        END
    END GCLK
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  24.85 5.40 26.35 6.30 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.55 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END CLK
    PIN CGOBS
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M2M ;
        RECT  18.50 2.70 19.10 8.45 ;
        RECT  18.50 2.70 19.30 3.80 ;
        RECT  18.50 7.35 19.30 8.45 ;
        LAYER M1M ;
        RECT  18.45 2.80 19.40 4.10 ;
        RECT  18.45 7.35 19.40 8.95 ;
        END
    END CGOBS
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.10 2.50 11.00 ;
        RECT  4.50 7.20 5.20 11.00 ;
        RECT  4.50 9.40 8.30 11.00 ;
        RECT  12.95 7.15 13.45 11.00 ;
        RECT  12.95 7.15 13.65 8.75 ;
        RECT  11.95 10.00 14.15 11.00 ;
        RECT  17.30 7.35 17.85 11.00 ;
        RECT  17.30 7.35 18.00 8.95 ;
        RECT  20.30 7.30 21.00 11.00 ;
        RECT  25.00 7.75 25.90 11.00 ;
        RECT  0.00 11.00 29.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.50 ;
        RECT  4.50 2.00 5.20 4.50 ;
        RECT  6.00 2.00 6.70 4.50 ;
        RECT  7.55 2.00 8.25 4.40 ;
        RECT  10.25 2.00 10.95 4.40 ;
        RECT  13.10 2.00 13.80 4.40 ;
        RECT  17.30 2.00 18.00 4.05 ;
        RECT  20.30 2.00 21.00 4.10 ;
        RECT  25.00 2.00 25.70 4.00 ;
        RECT  27.70 2.00 28.40 4.00 ;
        RECT  0.00 0.00 29.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.15 6.05 4.85 6.75 ;
        RECT  4.15 6.25 7.35 6.75 ;
        RECT  6.85 6.25 7.35 7.80 ;
        RECT  8.90 2.70 9.40 7.80 ;
        RECT  8.90 2.70 9.60 4.50 ;
        RECT  6.85 7.10 10.65 7.80 ;
        RECT  9.95 7.10 10.65 10.55 ;
        RECT  11.75 3.75 12.30 8.90 ;
        RECT  11.60 7.15 12.30 8.90 ;
        RECT  11.75 3.75 12.45 4.50 ;
        RECT  13.45 6.00 14.15 6.70 ;
        RECT  11.75 6.20 14.15 6.70 ;
        RECT  14.35 7.15 15.10 8.75 ;
        RECT  14.60 3.70 15.10 9.95 ;
        RECT  14.45 3.70 15.15 4.45 ;
        RECT  14.60 9.45 16.30 9.95 ;
        RECT  15.60 9.45 16.30 10.15 ;
        RECT  15.95 3.40 16.45 8.90 ;
        RECT  15.95 7.30 16.65 8.90 ;
        RECT  15.95 3.40 16.70 4.10 ;
        RECT  17.80 6.10 18.50 6.85 ;
        RECT  15.95 5.15 21.40 5.65 ;
        RECT  20.70 5.15 21.40 5.85 ;
        RECT  22.05 3.30 22.55 6.85 ;
        RECT  17.80 6.35 23.15 6.85 ;
        RECT  22.20 9.50 22.90 10.20 ;
        RECT  22.65 6.35 23.15 8.75 ;
        RECT  22.05 3.30 23.35 4.00 ;
        RECT  22.65 7.15 23.35 8.75 ;
        RECT  23.30 4.55 24.30 5.25 ;
        RECT  23.80 4.55 24.30 10.00 ;
        RECT  22.20 9.50 24.30 10.00 ;
        RECT  26.35 3.35 27.05 4.05 ;
        RECT  26.55 3.35 27.05 4.95 ;
        RECT  27.55 7.15 28.25 10.55 ;
        RECT  26.55 4.45 28.85 4.95 ;
        RECT  28.35 4.45 28.85 7.65 ;
        RECT  27.55 7.15 28.85 7.65 ;
        RECT  28.35 5.45 29.05 6.15 ;
        LAYER V1M ;
        RECT  18.40 6.65 19.40 7.65 ;
        RECT  18.40 7.95 19.40 8.95 ;
        RECT  18.40 2.75 19.40 3.75 ;
    END
END LSOGCNX8
MACRO LSOGCPX1
    CLASS CORE ;
    FOREIGN LSOGCPX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 26.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.45 3.35 1.15 4.15 ;
        RECT  0.25 5.35 1.15 6.35 ;
        RECT  0.65 3.35 1.15 8.75 ;
        RECT  0.45 7.10 1.15 8.75 ;
        END
    END GCLK
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END CLK
    PIN CGOBS
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  13.70 3.40 14.40 4.10 ;
        RECT  13.70 7.35 14.40 8.95 ;
        RECT  13.90 3.40 14.40 10.20 ;
        RECT  13.90 9.30 15.15 10.20 ;
        END
    END CGOBS
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  21.25 5.40 22.60 6.30 ;
        END
    END SE
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  15.30 8.30 16.10 8.85 ;
        RECT  1.80 7.25 2.50 11.00 ;
        RECT  4.65 7.15 5.35 11.00 ;
        RECT  3.45 9.05 5.35 11.00 ;
        RECT  7.60 7.15 8.10 11.00 ;
        RECT  7.60 7.15 8.30 8.75 ;
        RECT  0.85 10.10 8.65 11.00 ;
        RECT  12.35 7.35 12.90 11.00 ;
        RECT  12.35 7.35 13.05 8.95 ;
        RECT  15.60 7.25 16.00 11.00 ;
        RECT  15.30 7.25 16.00 8.85 ;
        RECT  15.60 8.30 16.10 11.00 ;
        RECT  20.00 7.75 20.90 11.00 ;
        RECT  24.05 7.15 24.75 11.00 ;
        RECT  0.00 11.00 26.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.10 ;
        RECT  8.10 2.00 8.80 4.40 ;
        RECT  12.35 2.00 13.05 4.05 ;
        RECT  15.30 2.00 16.00 4.10 ;
        RECT  20.00 2.00 20.70 4.00 ;
        RECT  22.70 2.00 23.40 4.00 ;
        RECT  0.00 0.00 26.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.60 6.05 2.30 6.75 ;
        RECT  1.60 6.20 3.90 6.75 ;
        RECT  3.40 4.45 3.90 7.85 ;
        RECT  3.30 6.20 3.90 7.85 ;
        RECT  3.30 7.15 4.00 7.85 ;
        RECT  4.30 3.40 5.00 4.95 ;
        RECT  3.40 4.45 5.00 4.95 ;
        RECT  6.40 6.20 6.95 8.90 ;
        RECT  6.75 3.75 6.95 8.90 ;
        RECT  6.25 7.15 6.95 8.90 ;
        RECT  6.75 3.75 7.30 6.70 ;
        RECT  6.75 3.75 7.45 4.50 ;
        RECT  8.00 6.00 8.70 6.70 ;
        RECT  6.40 6.20 8.70 6.70 ;
        RECT  9.00 7.15 9.75 8.75 ;
        RECT  9.25 3.70 9.75 10.55 ;
        RECT  9.15 7.15 9.75 10.55 ;
        RECT  9.15 9.85 9.85 10.55 ;
        RECT  9.25 3.70 10.15 4.45 ;
        RECT  11.00 3.40 11.50 8.90 ;
        RECT  11.00 3.40 11.70 4.10 ;
        RECT  11.00 7.30 11.70 8.90 ;
        RECT  11.00 5.30 13.40 5.80 ;
        RECT  12.70 5.30 13.40 6.00 ;
        RECT  14.95 6.10 15.65 6.80 ;
        RECT  17.05 3.30 17.55 6.80 ;
        RECT  14.95 6.30 18.15 6.80 ;
        RECT  17.20 9.50 17.90 10.20 ;
        RECT  17.65 6.30 18.15 8.75 ;
        RECT  17.05 3.30 18.35 4.00 ;
        RECT  17.65 7.15 18.35 8.75 ;
        RECT  18.30 4.55 19.30 5.25 ;
        RECT  18.80 4.55 19.30 10.00 ;
        RECT  17.20 9.50 19.30 10.00 ;
        RECT  21.35 3.35 22.05 4.05 ;
        RECT  21.55 3.35 22.05 4.95 ;
        RECT  21.55 4.45 23.60 4.95 ;
        RECT  23.10 4.45 23.25 10.55 ;
        RECT  22.55 7.15 23.25 10.55 ;
        RECT  23.10 4.45 23.60 7.65 ;
        RECT  22.55 7.15 23.60 7.65 ;
        RECT  23.10 5.45 23.85 6.15 ;
        RECT  24.05 3.30 24.75 4.00 ;
        RECT  25.40 3.30 25.90 8.95 ;
        RECT  25.30 3.30 26.00 4.00 ;
        RECT  24.05 3.50 26.00 4.00 ;
        RECT  25.40 7.20 26.10 8.95 ;
    END
END LSOGCPX1
MACRO LSOGCPX2
    CLASS CORE ;
    FOREIGN LSOGCPX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 26.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.50 1.15 4.45 ;
        RECT  0.25 5.35 1.15 6.35 ;
        RECT  0.65 2.50 1.15 10.55 ;
        RECT  0.45 7.10 1.15 10.55 ;
        END
    END GCLK
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END CLK
    PIN CGOBS
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  13.70 3.40 14.40 4.10 ;
        RECT  13.70 7.35 14.40 8.95 ;
        RECT  13.90 3.40 14.40 10.20 ;
        RECT  13.90 9.30 15.15 10.20 ;
        END
    END CGOBS
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  21.25 5.40 22.60 6.30 ;
        END
    END SE
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  15.30 8.30 16.10 8.85 ;
        RECT  1.80 7.25 2.50 11.00 ;
        RECT  4.65 7.15 5.35 11.00 ;
        RECT  3.45 9.05 5.35 11.00 ;
        RECT  7.60 7.15 8.10 11.00 ;
        RECT  7.60 7.15 8.30 8.75 ;
        RECT  3.45 10.10 8.65 11.00 ;
        RECT  12.35 7.35 12.90 11.00 ;
        RECT  12.35 7.35 13.05 8.95 ;
        RECT  15.60 7.25 16.00 11.00 ;
        RECT  15.30 7.25 16.00 8.85 ;
        RECT  15.60 8.30 16.10 11.00 ;
        RECT  20.00 7.75 20.90 11.00 ;
        RECT  24.05 7.15 24.75 11.00 ;
        RECT  0.00 11.00 26.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 3.90 ;
        RECT  8.10 2.00 8.80 4.40 ;
        RECT  12.35 2.00 13.05 4.05 ;
        RECT  15.30 2.00 16.00 4.10 ;
        RECT  20.00 2.00 20.70 4.00 ;
        RECT  22.70 2.00 23.40 4.00 ;
        RECT  0.00 0.00 26.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.60 6.05 2.30 6.75 ;
        RECT  1.60 6.20 3.90 6.75 ;
        RECT  3.40 4.45 3.90 7.85 ;
        RECT  3.30 6.20 3.90 7.85 ;
        RECT  3.30 7.15 4.00 7.85 ;
        RECT  4.30 3.40 5.00 4.95 ;
        RECT  3.40 4.45 5.00 4.95 ;
        RECT  6.40 6.20 6.95 8.90 ;
        RECT  6.75 3.75 6.95 8.90 ;
        RECT  6.25 7.15 6.95 8.90 ;
        RECT  6.75 3.75 7.30 6.70 ;
        RECT  6.75 3.75 7.45 4.50 ;
        RECT  8.00 6.00 8.70 6.70 ;
        RECT  6.40 6.20 8.70 6.70 ;
        RECT  9.00 7.15 9.75 8.75 ;
        RECT  9.25 3.70 9.75 10.55 ;
        RECT  9.15 7.15 9.75 10.55 ;
        RECT  9.15 9.85 9.85 10.55 ;
        RECT  9.25 3.70 10.15 4.45 ;
        RECT  11.00 3.40 11.50 8.90 ;
        RECT  11.00 3.40 11.70 4.10 ;
        RECT  11.00 7.30 11.70 8.90 ;
        RECT  11.00 5.30 13.40 5.80 ;
        RECT  12.70 5.30 13.40 6.00 ;
        RECT  14.95 6.10 15.65 6.80 ;
        RECT  17.05 3.30 17.55 6.80 ;
        RECT  14.95 6.30 18.15 6.80 ;
        RECT  17.20 9.50 17.90 10.20 ;
        RECT  17.65 6.30 18.15 8.75 ;
        RECT  17.05 3.30 18.35 4.00 ;
        RECT  17.65 7.15 18.35 8.75 ;
        RECT  18.30 4.55 19.30 5.25 ;
        RECT  18.80 4.55 19.30 10.00 ;
        RECT  17.20 9.50 19.30 10.00 ;
        RECT  21.35 3.35 22.05 4.05 ;
        RECT  21.55 3.35 22.05 4.95 ;
        RECT  21.55 4.45 23.60 4.95 ;
        RECT  23.10 4.45 23.25 10.55 ;
        RECT  22.55 7.15 23.25 10.55 ;
        RECT  23.10 4.45 23.60 7.65 ;
        RECT  22.55 7.15 23.60 7.65 ;
        RECT  23.10 5.45 23.85 6.15 ;
        RECT  24.05 3.30 24.75 4.00 ;
        RECT  25.40 3.30 25.90 8.95 ;
        RECT  25.30 3.30 26.00 4.00 ;
        RECT  24.05 3.50 26.00 4.00 ;
        RECT  25.40 7.20 26.10 8.95 ;
    END
END LSOGCPX2
MACRO LSOGCPX3
    CLASS CORE ;
    FOREIGN LSOGCPX3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 28.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.35 1.15 6.35 ;
        RECT  0.25 5.65 2.45 6.15 ;
        RECT  1.95 4.45 2.45 9.40 ;
        RECT  1.95 7.10 2.65 9.40 ;
        RECT  2.50 3.15 3.00 4.95 ;
        RECT  1.95 4.45 3.00 4.95 ;
        RECT  2.50 3.15 3.20 3.85 ;
        END
    END GCLK
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  21.25 5.40 22.15 6.30 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END CLK
    PIN CGOBS
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  15.10 3.40 15.80 4.10 ;
        RECT  15.10 7.35 15.80 8.95 ;
        RECT  15.30 3.40 15.80 10.20 ;
        RECT  15.30 9.30 16.55 10.20 ;
        END
    END CGOBS
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  22.65 5.40 24.00 6.30 ;
        END
    END SE
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  16.70 8.30 17.50 8.85 ;
        RECT  0.60 7.10 1.30 11.00 ;
        RECT  3.30 7.25 4.00 11.00 ;
        RECT  6.15 7.15 6.85 11.00 ;
        RECT  9.00 7.15 9.50 11.00 ;
        RECT  9.00 7.15 9.70 8.75 ;
        RECT  4.85 10.10 10.05 11.00 ;
        RECT  13.75 7.35 14.30 11.00 ;
        RECT  13.75 7.35 14.45 8.95 ;
        RECT  17.00 7.25 17.40 11.00 ;
        RECT  16.70 7.25 17.40 8.85 ;
        RECT  17.00 8.30 17.50 11.00 ;
        RECT  21.40 7.75 22.30 11.00 ;
        RECT  25.45 7.15 26.15 11.00 ;
        RECT  0.00 11.00 28.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.15 2.00 1.85 3.85 ;
        RECT  4.00 2.00 4.70 4.00 ;
        RECT  9.50 2.00 10.20 4.40 ;
        RECT  13.75 2.00 14.45 4.05 ;
        RECT  16.70 2.00 17.40 4.10 ;
        RECT  21.40 2.00 22.10 4.00 ;
        RECT  24.10 2.00 24.80 4.00 ;
        RECT  0.00 0.00 28.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.10 6.05 3.80 6.75 ;
        RECT  3.10 6.20 5.30 6.75 ;
        RECT  4.80 4.45 5.30 8.75 ;
        RECT  4.80 7.15 5.50 8.75 ;
        RECT  6.35 2.55 7.05 4.95 ;
        RECT  4.80 4.45 7.05 4.95 ;
        RECT  7.80 6.20 8.35 8.90 ;
        RECT  8.15 3.75 8.35 8.90 ;
        RECT  7.65 7.15 8.35 8.90 ;
        RECT  8.15 3.75 8.70 6.70 ;
        RECT  8.15 3.75 8.85 4.50 ;
        RECT  9.40 6.00 10.10 6.70 ;
        RECT  7.80 6.20 10.10 6.70 ;
        RECT  10.40 7.15 11.15 8.75 ;
        RECT  10.65 3.70 11.15 10.55 ;
        RECT  10.55 7.15 11.15 10.55 ;
        RECT  10.55 9.85 11.25 10.55 ;
        RECT  10.65 3.70 11.55 4.45 ;
        RECT  12.40 3.40 12.90 8.90 ;
        RECT  12.40 3.40 13.10 4.10 ;
        RECT  12.40 7.30 13.10 8.90 ;
        RECT  12.40 5.30 14.80 5.80 ;
        RECT  14.10 5.30 14.80 6.00 ;
        RECT  16.35 6.10 17.05 6.80 ;
        RECT  18.45 3.30 18.95 6.80 ;
        RECT  16.35 6.30 19.55 6.80 ;
        RECT  18.60 9.50 19.30 10.20 ;
        RECT  19.05 6.30 19.55 8.75 ;
        RECT  18.45 3.30 19.75 4.00 ;
        RECT  19.05 7.15 19.75 8.75 ;
        RECT  19.70 4.55 20.70 5.25 ;
        RECT  20.20 4.55 20.70 10.00 ;
        RECT  18.60 9.50 20.70 10.00 ;
        RECT  22.75 3.35 23.45 4.05 ;
        RECT  22.95 3.35 23.45 4.95 ;
        RECT  22.95 4.45 25.00 4.95 ;
        RECT  24.50 4.45 24.65 10.55 ;
        RECT  23.95 7.15 24.65 10.55 ;
        RECT  24.50 4.45 25.00 7.65 ;
        RECT  23.95 7.15 25.00 7.65 ;
        RECT  24.50 5.45 25.25 6.15 ;
        RECT  25.45 3.30 26.15 4.00 ;
        RECT  26.80 3.30 27.30 8.95 ;
        RECT  26.70 3.30 27.40 4.00 ;
        RECT  25.45 3.50 27.40 4.00 ;
        RECT  26.80 7.20 27.50 8.95 ;
    END
END LSOGCPX3
MACRO LSOGCPX4
    CLASS CORE ;
    FOREIGN LSOGCPX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 28.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.35 1.15 6.35 ;
        RECT  0.25 5.65 2.45 6.15 ;
        RECT  1.95 4.45 2.45 10.55 ;
        RECT  1.95 7.10 2.65 10.55 ;
        RECT  2.65 2.55 3.15 4.95 ;
        RECT  1.95 4.45 3.15 4.95 ;
        RECT  2.65 2.55 3.35 4.55 ;
        RECT  1.95 4.45 3.35 4.55 ;
        END
    END GCLK
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  21.25 5.40 22.15 6.30 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END CLK
    PIN CGOBS
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  15.10 3.40 15.80 4.10 ;
        RECT  15.10 7.35 15.80 8.95 ;
        RECT  15.30 3.40 15.80 10.20 ;
        RECT  15.30 9.30 16.55 10.20 ;
        END
    END CGOBS
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  22.65 5.40 24.00 6.30 ;
        END
    END SE
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  16.70 8.30 17.50 8.85 ;
        RECT  0.60 7.10 1.30 11.00 ;
        RECT  3.30 7.25 4.00 11.00 ;
        RECT  6.15 7.15 6.85 11.00 ;
        RECT  9.00 7.15 9.50 11.00 ;
        RECT  9.00 7.15 9.70 8.75 ;
        RECT  4.85 10.10 10.05 11.00 ;
        RECT  13.75 7.35 14.30 11.00 ;
        RECT  13.75 7.35 14.45 8.95 ;
        RECT  17.00 7.25 17.40 11.00 ;
        RECT  16.70 7.25 17.40 8.85 ;
        RECT  17.00 8.30 17.50 11.00 ;
        RECT  21.40 7.75 22.30 11.00 ;
        RECT  25.45 7.15 26.15 11.00 ;
        RECT  0.00 11.00 28.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.30 2.00 2.00 4.00 ;
        RECT  4.00 2.00 4.70 4.00 ;
        RECT  9.50 2.00 10.20 4.40 ;
        RECT  13.75 2.00 14.45 4.05 ;
        RECT  16.70 2.00 17.40 4.10 ;
        RECT  21.40 2.00 22.10 4.00 ;
        RECT  24.10 2.00 24.80 4.00 ;
        RECT  0.00 0.00 28.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.10 6.05 3.80 6.75 ;
        RECT  3.10 6.20 5.30 6.75 ;
        RECT  4.80 4.45 5.30 8.75 ;
        RECT  4.80 7.15 5.50 8.75 ;
        RECT  6.35 2.55 7.05 4.95 ;
        RECT  4.80 4.45 7.05 4.95 ;
        RECT  7.80 6.20 8.35 8.90 ;
        RECT  8.15 3.75 8.35 8.90 ;
        RECT  7.65 7.15 8.35 8.90 ;
        RECT  8.15 3.75 8.70 6.70 ;
        RECT  8.15 3.75 8.85 4.50 ;
        RECT  9.40 6.00 10.10 6.70 ;
        RECT  7.80 6.20 10.10 6.70 ;
        RECT  10.40 7.15 11.15 8.75 ;
        RECT  10.65 3.70 11.15 10.55 ;
        RECT  10.55 7.15 11.15 10.55 ;
        RECT  10.55 9.85 11.25 10.55 ;
        RECT  10.65 3.70 11.55 4.45 ;
        RECT  12.40 3.40 12.90 8.90 ;
        RECT  12.40 3.40 13.10 4.10 ;
        RECT  12.40 7.30 13.10 8.90 ;
        RECT  12.40 5.30 14.80 5.80 ;
        RECT  14.10 5.30 14.80 6.00 ;
        RECT  16.35 6.10 17.05 6.80 ;
        RECT  18.45 3.30 18.95 6.80 ;
        RECT  16.35 6.30 19.55 6.80 ;
        RECT  18.60 9.50 19.30 10.20 ;
        RECT  19.05 6.30 19.55 8.75 ;
        RECT  18.45 3.30 19.75 4.00 ;
        RECT  19.05 7.15 19.75 8.75 ;
        RECT  19.70 4.55 20.70 5.25 ;
        RECT  20.20 4.55 20.70 10.00 ;
        RECT  18.60 9.50 20.70 10.00 ;
        RECT  22.75 3.35 23.45 4.05 ;
        RECT  22.95 3.35 23.45 4.95 ;
        RECT  22.95 4.45 25.00 4.95 ;
        RECT  24.50 4.45 24.65 10.55 ;
        RECT  23.95 7.15 24.65 10.55 ;
        RECT  24.50 4.45 25.00 7.65 ;
        RECT  23.95 7.15 25.00 7.65 ;
        RECT  24.50 5.45 25.25 6.15 ;
        RECT  25.45 3.30 26.15 4.00 ;
        RECT  26.80 3.30 27.30 8.95 ;
        RECT  26.70 3.30 27.40 4.00 ;
        RECT  25.45 3.50 27.40 4.00 ;
        RECT  26.80 7.20 27.50 8.95 ;
    END
END LSOGCPX4
MACRO LSOGCPX8
    CLASS CORE ;
    FOREIGN LSOGCPX8 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 29.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.50 1.20 4.55 ;
        RECT  1.00 2.50 1.20 10.55 ;
        RECT  0.70 2.50 1.20 6.10 ;
        RECT  1.00 5.60 1.50 10.55 ;
        RECT  0.80 7.10 1.50 10.55 ;
        RECT  1.65 5.35 2.55 6.35 ;
        RECT  1.00 5.60 2.55 6.35 ;
        RECT  3.15 2.50 3.70 6.60 ;
        RECT  3.15 6.10 4.00 6.60 ;
        RECT  3.50 2.50 3.70 10.55 ;
        RECT  0.70 5.60 3.70 6.10 ;
        RECT  3.15 2.50 3.85 4.50 ;
        RECT  3.50 6.10 4.00 10.55 ;
        RECT  3.50 7.10 4.20 10.55 ;
        END
    END GCLK
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  22.65 5.40 23.55 6.30 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.85 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END CLK
    PIN CGOBS
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  16.50 3.40 17.20 4.10 ;
        RECT  16.50 7.35 17.20 8.95 ;
        RECT  16.70 3.40 17.20 10.20 ;
        RECT  16.70 9.30 17.95 10.20 ;
        END
    END CGOBS
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  24.05 5.40 25.40 6.30 ;
        END
    END SE
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  18.10 8.30 18.90 8.85 ;
        RECT  2.15 7.10 2.85 11.00 ;
        RECT  4.85 7.25 5.55 11.00 ;
        RECT  7.55 7.35 8.25 11.00 ;
        RECT  10.40 7.15 10.90 11.00 ;
        RECT  10.40 7.15 11.10 8.75 ;
        RECT  9.40 10.00 11.45 11.00 ;
        RECT  15.15 7.35 15.70 11.00 ;
        RECT  15.15 7.35 15.85 8.95 ;
        RECT  18.40 7.25 18.80 11.00 ;
        RECT  18.10 7.25 18.80 8.85 ;
        RECT  18.40 8.30 18.90 11.00 ;
        RECT  22.80 7.75 23.70 11.00 ;
        RECT  26.85 7.15 27.55 11.00 ;
        RECT  0.00 11.00 29.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.50 ;
        RECT  4.50 2.00 5.20 4.50 ;
        RECT  10.90 2.00 11.60 4.40 ;
        RECT  15.15 2.00 15.85 4.05 ;
        RECT  18.10 2.00 18.80 4.10 ;
        RECT  22.80 2.00 23.50 4.00 ;
        RECT  25.50 2.00 26.20 4.00 ;
        RECT  0.00 0.00 29.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.15 4.95 4.85 5.65 ;
        RECT  4.15 5.10 6.70 5.65 ;
        RECT  6.20 3.80 6.70 10.55 ;
        RECT  6.20 8.05 6.90 10.55 ;
        RECT  8.00 2.50 8.75 4.50 ;
        RECT  6.20 3.80 8.75 4.50 ;
        RECT  9.20 6.20 9.75 8.90 ;
        RECT  9.55 3.75 9.75 8.90 ;
        RECT  9.05 7.15 9.75 8.90 ;
        RECT  9.55 3.75 10.10 6.70 ;
        RECT  9.55 3.75 10.25 4.50 ;
        RECT  10.80 6.00 11.50 6.70 ;
        RECT  9.20 6.20 11.50 6.70 ;
        RECT  11.80 7.15 12.55 8.75 ;
        RECT  12.05 3.70 12.55 10.55 ;
        RECT  11.95 7.15 12.55 10.55 ;
        RECT  11.95 9.85 12.65 10.55 ;
        RECT  12.05 3.70 12.95 4.45 ;
        RECT  13.80 3.40 14.30 8.90 ;
        RECT  13.80 3.40 14.50 4.10 ;
        RECT  13.80 7.30 14.50 8.90 ;
        RECT  13.80 5.30 16.20 5.80 ;
        RECT  15.50 5.30 16.20 6.00 ;
        RECT  17.75 6.10 18.45 6.80 ;
        RECT  19.85 3.30 20.35 6.80 ;
        RECT  17.75 6.30 20.95 6.80 ;
        RECT  20.00 9.50 20.70 10.20 ;
        RECT  20.45 6.30 20.95 8.75 ;
        RECT  19.85 3.30 21.15 4.00 ;
        RECT  20.45 7.15 21.15 8.75 ;
        RECT  21.10 4.55 22.10 5.25 ;
        RECT  21.60 4.55 22.10 10.00 ;
        RECT  20.00 9.50 22.10 10.00 ;
        RECT  24.15 3.35 24.85 4.05 ;
        RECT  24.35 3.35 24.85 4.95 ;
        RECT  24.35 4.45 26.40 4.95 ;
        RECT  25.90 4.45 26.05 10.55 ;
        RECT  25.35 7.15 26.05 10.55 ;
        RECT  25.90 4.45 26.40 7.65 ;
        RECT  25.35 7.15 26.40 7.65 ;
        RECT  25.90 5.45 26.65 6.15 ;
        RECT  26.85 3.30 27.55 4.00 ;
        RECT  28.20 3.30 28.70 8.95 ;
        RECT  28.10 3.30 28.80 4.00 ;
        RECT  26.85 3.50 28.80 4.00 ;
        RECT  28.20 7.20 28.90 8.95 ;
    END
END LSOGCPX8
MACRO MU2IX1
    CLASS CORE ;
    FOREIGN MU2IX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN S
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END S
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.85 2.80 6.05 4.45 ;
        RECT  4.85 7.70 5.55 10.55 ;
        RECT  5.55 2.80 6.05 8.20 ;
        RECT  4.85 7.70 6.05 8.20 ;
        RECT  4.85 2.80 6.75 3.70 ;
        END
    END Q
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END IN1
    PIN IN0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END IN0
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.55 10.10 1.25 11.00 ;
        RECT  2.50 7.70 3.20 11.00 ;
        RECT  7.20 7.30 7.90 11.00 ;
        RECT  0.00 11.00 8.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.50 2.00 3.20 4.40 ;
        RECT  7.20 2.00 7.90 4.40 ;
        RECT  0.00 0.00 8.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.00 3.75 1.20 8.80 ;
        RECT  0.70 3.75 1.20 7.25 ;
        RECT  0.70 3.75 1.70 4.50 ;
        RECT  1.00 6.75 1.70 8.80 ;
        RECT  4.40 5.40 4.90 7.25 ;
        RECT  0.70 6.75 4.90 7.25 ;
        RECT  4.40 5.40 5.10 6.10 ;
    END
END MU2IX1
MACRO MU2IX2
    CLASS CORE ;
    FOREIGN MU2IX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN S
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.25 ;
        PORT
        LAYER M1M ;
        RECT  1.50 5.40 2.55 6.30 ;
        END
    END S
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  6.05 2.45 6.75 3.90 ;
        RECT  6.05 8.70 6.75 10.55 ;
        RECT  8.75 2.45 9.45 4.50 ;
        RECT  8.95 2.45 9.45 10.55 ;
        RECT  8.75 7.70 9.45 10.55 ;
        RECT  8.65 5.40 9.55 6.30 ;
        RECT  6.05 2.45 12.15 2.95 ;
        RECT  11.45 2.45 12.15 3.90 ;
        RECT  11.45 7.75 12.15 10.55 ;
        RECT  6.05 10.05 12.15 10.55 ;
        END
    END Q
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.20 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END IN1
    PIN IN0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.20 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END IN0
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 7.70 2.55 11.00 ;
        RECT  4.55 8.65 5.25 11.00 ;
        RECT  12.95 7.75 13.65 11.00 ;
        RECT  15.65 7.30 16.35 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 2.00 2.55 4.40 ;
        RECT  4.55 2.00 5.25 3.90 ;
        RECT  12.95 2.00 13.65 3.90 ;
        RECT  15.65 2.00 16.35 4.40 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.75 0.95 8.80 ;
        RECT  0.45 3.75 1.15 4.50 ;
        RECT  0.45 6.75 1.15 8.80 ;
        RECT  3.20 2.70 3.90 4.90 ;
        RECT  3.20 7.70 3.90 10.55 ;
        RECT  4.95 5.40 5.45 7.25 ;
        RECT  0.45 6.75 5.45 7.25 ;
        RECT  4.95 5.40 5.65 6.10 ;
        RECT  3.20 7.70 8.10 8.20 ;
        RECT  7.40 3.45 8.10 4.90 ;
        RECT  3.20 4.40 8.10 4.90 ;
        RECT  7.40 7.70 8.10 9.60 ;
        RECT  10.10 3.45 10.80 4.90 ;
        RECT  10.10 6.80 10.80 9.60 ;
        RECT  10.10 6.80 15.00 7.30 ;
        RECT  14.30 2.70 15.00 4.90 ;
        RECT  10.10 4.40 15.00 4.90 ;
        RECT  14.30 6.80 15.00 10.55 ;
    END
END MU2IX2
MACRO MU2IX4
    CLASS CORE ;
    FOREIGN MU2IX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 28.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN S
        DIRECTION INPUT ;
        ANTENNAGATEAREA 10.50 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END S
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  9.05 2.45 9.75 3.90 ;
        RECT  9.05 7.55 9.75 10.55 ;
        RECT  11.75 2.45 12.45 4.50 ;
        RECT  11.75 7.55 12.45 10.55 ;
        RECT  14.25 5.40 15.15 6.30 ;
        RECT  14.45 2.45 15.15 10.55 ;
        RECT  17.15 2.45 17.85 4.50 ;
        RECT  17.15 7.55 17.85 10.55 ;
        RECT  9.05 2.45 20.55 2.95 ;
        RECT  19.85 2.45 20.55 4.50 ;
        RECT  19.85 7.55 20.55 10.55 ;
        RECT  9.05 10.05 20.55 10.55 ;
        END
    END Q
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 8.40 ;
        PORT
        LAYER M1M ;
        RECT  25.45 5.40 26.35 6.30 ;
        END
    END IN1
    PIN IN0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 8.40 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END IN0
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.15 7.70 2.85 11.00 ;
        RECT  4.85 8.65 5.55 11.00 ;
        RECT  7.55 7.55 8.25 11.00 ;
        RECT  21.35 7.50 22.05 11.00 ;
        RECT  24.05 7.75 24.75 11.00 ;
        RECT  26.75 7.30 27.45 11.00 ;
        RECT  0.00 11.00 28.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.15 2.00 2.85 4.40 ;
        RECT  4.85 2.00 5.55 3.90 ;
        RECT  7.55 2.00 8.25 3.90 ;
        RECT  21.35 2.00 22.05 4.50 ;
        RECT  24.05 2.00 24.75 3.90 ;
        RECT  26.75 2.00 27.45 4.40 ;
        RECT  0.00 0.00 28.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.65 2.75 1.15 10.50 ;
        RECT  0.65 2.75 1.35 4.50 ;
        RECT  0.65 6.75 1.35 10.50 ;
        RECT  3.50 2.70 4.20 4.90 ;
        RECT  3.50 7.70 4.20 10.55 ;
        RECT  4.70 5.60 5.20 7.25 ;
        RECT  0.65 6.75 5.20 7.25 ;
        RECT  3.50 7.70 6.90 8.20 ;
        RECT  6.20 2.70 6.90 4.90 ;
        RECT  6.20 6.55 6.90 10.55 ;
        RECT  9.25 5.40 9.95 6.10 ;
        RECT  4.70 5.60 9.95 6.10 ;
        RECT  3.50 4.40 11.10 4.90 ;
        RECT  10.40 3.45 11.10 5.50 ;
        RECT  10.40 6.55 11.10 9.60 ;
        RECT  6.20 6.55 13.80 7.05 ;
        RECT  13.10 3.45 13.80 5.50 ;
        RECT  10.40 5.00 13.80 5.50 ;
        RECT  13.10 6.55 13.80 9.60 ;
        RECT  15.80 3.45 16.50 5.50 ;
        RECT  15.80 6.55 16.50 9.60 ;
        RECT  18.50 3.45 19.20 5.50 ;
        RECT  18.50 6.55 19.20 9.60 ;
        RECT  15.80 6.55 23.40 7.05 ;
        RECT  15.80 6.80 26.10 7.05 ;
        RECT  22.70 2.70 23.40 5.50 ;
        RECT  15.80 5.00 23.40 5.50 ;
        RECT  22.70 6.55 23.40 10.55 ;
        RECT  22.70 6.80 26.10 7.30 ;
        RECT  25.40 2.70 26.10 4.90 ;
        RECT  22.70 4.40 26.10 4.90 ;
        RECT  25.40 6.80 26.10 10.55 ;
    END
END MU2IX4
MACRO MU2X1
    CLASS CORE ;
    FOREIGN MU2X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN S
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END S
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.20 3.00 8.90 3.75 ;
        RECT  8.40 3.00 8.90 9.70 ;
        RECT  8.20 8.10 8.90 9.70 ;
        RECT  8.40 5.40 9.55 6.30 ;
        END
    END Q
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END IN1
    PIN IN0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END IN0
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.15 8.05 2.85 11.00 ;
        RECT  6.85 8.15 7.55 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.15 2.00 2.85 3.75 ;
        RECT  6.85 2.00 7.55 3.75 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.70 3.05 1.20 9.65 ;
        RECT  0.70 3.05 1.50 4.75 ;
        RECT  0.70 8.05 1.50 9.65 ;
        RECT  0.70 4.25 4.75 4.75 ;
        RECT  4.05 4.25 4.75 4.95 ;
        RECT  4.50 3.05 5.70 3.75 ;
        RECT  4.50 7.20 5.20 9.65 ;
        RECT  5.20 3.05 5.70 4.75 ;
        RECT  5.20 4.25 7.70 4.75 ;
        RECT  7.20 4.25 7.70 7.70 ;
        RECT  4.50 7.20 7.70 7.70 ;
        RECT  7.20 5.50 7.95 6.20 ;
    END
END MU2X1
MACRO MU2X2
    CLASS CORE ;
    FOREIGN MU2X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN S
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END S
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.35 2.45 9.05 4.05 ;
        RECT  8.55 2.45 9.05 10.50 ;
        RECT  8.35 7.10 9.05 10.50 ;
        RECT  8.55 5.40 9.55 6.30 ;
        END
    END Q
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END IN1
    PIN IN0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END IN0
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.15 8.05 2.85 11.00 ;
        RECT  7.00 7.70 7.70 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.15 2.00 2.85 3.75 ;
        RECT  7.00 2.00 7.70 4.00 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.70 3.05 1.20 9.65 ;
        RECT  0.70 3.05 1.50 4.75 ;
        RECT  0.70 8.05 1.50 9.65 ;
        RECT  0.70 4.25 4.75 4.75 ;
        RECT  4.05 4.25 4.75 4.95 ;
        RECT  4.50 3.05 5.70 3.75 ;
        RECT  4.50 6.75 5.20 9.65 ;
        RECT  5.20 3.05 5.70 4.95 ;
        RECT  5.20 4.45 7.70 4.95 ;
        RECT  7.20 4.45 7.70 7.25 ;
        RECT  4.50 6.75 7.70 7.25 ;
        RECT  7.20 5.50 7.95 6.20 ;
    END
END MU2X2
MACRO MU2X4
    CLASS CORE ;
    FOREIGN MU2X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN S
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END S
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.35 2.45 9.05 4.05 ;
        RECT  8.55 2.45 9.05 10.50 ;
        RECT  8.35 7.10 9.05 10.50 ;
        RECT  8.55 5.40 9.55 6.30 ;
        END
    END Q
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END IN1
    PIN IN0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END IN0
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.15 8.05 2.85 11.00 ;
        RECT  7.00 7.70 7.70 11.00 ;
        RECT  9.70 7.10 10.40 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.15 2.00 2.85 3.75 ;
        RECT  7.00 2.00 7.70 4.00 ;
        RECT  9.70 2.00 10.40 4.00 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.70 3.05 1.20 9.65 ;
        RECT  0.70 3.05 1.50 4.75 ;
        RECT  0.70 8.05 1.50 9.65 ;
        RECT  0.70 4.25 4.75 4.75 ;
        RECT  4.05 4.25 4.75 4.95 ;
        RECT  4.50 3.05 5.70 3.75 ;
        RECT  4.50 6.75 5.20 9.65 ;
        RECT  5.20 3.05 5.70 4.95 ;
        RECT  5.20 4.45 7.70 4.95 ;
        RECT  7.20 4.45 7.70 7.25 ;
        RECT  4.50 6.75 7.70 7.25 ;
        RECT  7.20 5.50 7.95 6.20 ;
    END
END MU2X4
MACRO MU4IX1
    CLASS CORE ;
    FOREIGN MU4IX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN S1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  17.05 6.70 17.95 7.60 ;
        RECT  16.85 6.90 17.95 7.60 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  0.25 6.70 1.15 7.60 ;
        END
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  21.20 3.75 21.90 4.50 ;
        RECT  21.40 3.75 21.90 8.90 ;
        RECT  21.20 7.10 21.90 8.90 ;
        RECT  21.25 5.40 22.15 6.30 ;
        END
    END Q
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.20 6.70 8.15 7.60 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  10.05 6.70 11.30 7.60 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 6.70 6.75 7.60 ;
        END
    END IN1
    PIN IN0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END IN0
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 9.10 2.55 11.00 ;
        RECT  6.55 8.50 7.25 11.00 ;
        RECT  11.25 8.40 11.95 11.00 ;
        RECT  15.95 8.45 16.65 11.00 ;
        RECT  19.85 7.10 20.55 11.00 ;
        RECT  18.80 10.10 21.95 11.00 ;
        RECT  0.00 11.00 22.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 2.00 2.55 4.15 ;
        RECT  6.55 2.00 7.25 4.15 ;
        RECT  11.25 2.00 11.95 4.15 ;
        RECT  15.95 2.00 16.65 4.20 ;
        RECT  19.85 2.00 20.55 4.50 ;
        RECT  0.00 0.00 22.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.50 3.55 1.20 5.50 ;
        RECT  0.50 8.15 1.20 10.25 ;
        RECT  1.70 5.00 2.20 8.65 ;
        RECT  0.50 8.15 2.20 8.65 ;
        RECT  0.50 5.00 4.45 5.50 ;
        RECT  3.75 5.00 4.45 5.70 ;
        RECT  4.20 3.55 5.40 4.25 ;
        RECT  4.20 8.65 4.90 10.25 ;
        RECT  4.90 3.55 5.40 9.15 ;
        RECT  4.20 8.65 5.40 9.15 ;
        RECT  7.75 2.55 8.25 5.10 ;
        RECT  4.90 4.60 8.25 5.10 ;
        RECT  8.90 3.55 9.60 4.25 ;
        RECT  9.10 3.55 9.60 10.00 ;
        RECT  8.90 8.40 9.60 10.00 ;
        RECT  7.75 2.55 10.70 3.05 ;
        RECT  10.20 2.55 10.70 5.10 ;
        RECT  10.20 4.60 12.40 5.10 ;
        RECT  11.70 4.60 12.40 5.30 ;
        RECT  13.60 3.55 14.30 5.25 ;
        RECT  13.60 7.40 14.30 10.05 ;
        RECT  9.10 5.75 15.40 6.25 ;
        RECT  14.70 5.75 15.40 6.45 ;
        RECT  13.60 4.75 16.40 5.25 ;
        RECT  15.90 4.75 16.40 7.90 ;
        RECT  13.60 7.40 16.40 7.90 ;
        RECT  17.30 8.30 18.00 10.05 ;
        RECT  17.70 5.55 18.40 6.25 ;
        RECT  15.90 5.75 18.40 6.25 ;
        RECT  17.30 3.55 19.35 4.25 ;
        RECT  18.85 3.55 19.35 8.80 ;
        RECT  17.30 8.30 19.35 8.80 ;
    END
END MU4IX1
MACRO MU4IX2
    CLASS CORE ;
    FOREIGN MU4IX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN S1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  17.05 6.70 17.95 7.60 ;
        RECT  16.85 6.90 17.95 7.60 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  0.25 6.70 1.15 7.60 ;
        END
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  21.20 2.70 21.90 4.50 ;
        RECT  21.40 2.70 21.90 10.50 ;
        RECT  21.20 7.10 21.90 10.50 ;
        RECT  21.25 5.40 22.15 6.30 ;
        END
    END Q
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.20 6.70 8.15 7.60 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  10.05 6.70 11.30 7.60 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 6.70 6.75 7.60 ;
        END
    END IN1
    PIN IN0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END IN0
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 9.10 2.55 11.00 ;
        RECT  6.55 8.50 7.25 11.00 ;
        RECT  11.25 8.40 11.95 11.00 ;
        RECT  15.95 8.45 16.65 11.00 ;
        RECT  19.85 7.10 20.55 11.00 ;
        RECT  0.00 11.00 22.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 2.00 2.55 4.15 ;
        RECT  6.55 2.00 7.25 4.15 ;
        RECT  11.25 2.00 11.95 4.15 ;
        RECT  15.95 2.00 16.65 4.20 ;
        RECT  19.85 2.00 20.55 4.50 ;
        RECT  0.00 0.00 22.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.50 3.55 1.20 5.50 ;
        RECT  0.50 8.15 1.20 10.25 ;
        RECT  1.70 5.00 2.20 8.65 ;
        RECT  0.50 8.15 2.20 8.65 ;
        RECT  0.50 5.00 4.45 5.50 ;
        RECT  3.75 5.00 4.45 5.70 ;
        RECT  4.20 3.55 5.40 4.25 ;
        RECT  4.20 8.65 4.90 10.25 ;
        RECT  4.90 3.55 5.40 9.15 ;
        RECT  4.20 8.65 5.40 9.15 ;
        RECT  7.75 2.55 8.25 5.10 ;
        RECT  4.90 4.60 8.25 5.10 ;
        RECT  8.90 3.55 9.60 4.25 ;
        RECT  9.10 3.55 9.60 10.00 ;
        RECT  8.90 8.40 9.60 10.00 ;
        RECT  7.75 2.55 10.70 3.05 ;
        RECT  10.20 2.55 10.70 5.10 ;
        RECT  10.20 4.60 12.40 5.10 ;
        RECT  11.70 4.60 12.40 5.30 ;
        RECT  13.60 3.55 14.30 5.25 ;
        RECT  13.60 7.40 14.30 10.05 ;
        RECT  9.10 5.75 15.40 6.25 ;
        RECT  14.70 5.75 15.40 6.45 ;
        RECT  13.60 4.75 16.40 5.25 ;
        RECT  15.90 4.75 16.40 7.90 ;
        RECT  13.60 7.40 16.40 7.90 ;
        RECT  17.30 8.30 18.00 10.05 ;
        RECT  17.70 5.55 18.40 6.25 ;
        RECT  15.90 5.75 18.40 6.25 ;
        RECT  17.30 3.55 19.35 4.25 ;
        RECT  18.85 3.55 19.35 8.80 ;
        RECT  17.30 8.30 19.35 8.80 ;
    END
END MU4IX2
MACRO MU4IX4
    CLASS CORE ;
    FOREIGN MU4IX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN S1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  17.05 6.70 17.95 7.60 ;
        RECT  16.85 6.90 17.95 7.60 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  0.25 6.70 1.15 7.60 ;
        END
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  21.20 2.70 21.90 4.50 ;
        RECT  21.40 2.70 21.90 10.50 ;
        RECT  21.20 7.10 21.90 10.50 ;
        RECT  21.25 5.40 22.15 6.30 ;
        END
    END Q
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.20 6.70 8.15 7.60 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  10.05 6.70 11.30 7.60 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 6.70 6.75 7.60 ;
        END
    END IN1
    PIN IN0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END IN0
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 9.10 2.55 11.00 ;
        RECT  6.55 8.50 7.25 11.00 ;
        RECT  11.25 8.40 11.95 11.00 ;
        RECT  15.95 8.45 16.65 11.00 ;
        RECT  19.85 7.10 20.55 11.00 ;
        RECT  22.55 7.10 23.25 11.00 ;
        RECT  0.00 11.00 23.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 2.00 2.55 4.15 ;
        RECT  6.55 2.00 7.25 4.15 ;
        RECT  11.25 2.00 11.95 4.15 ;
        RECT  15.95 2.00 16.65 4.20 ;
        RECT  19.85 2.00 20.55 4.50 ;
        RECT  22.55 2.00 23.25 4.50 ;
        RECT  0.00 0.00 23.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.50 3.55 1.20 5.50 ;
        RECT  0.50 8.15 1.20 10.25 ;
        RECT  1.70 5.00 2.20 8.65 ;
        RECT  0.50 8.15 2.20 8.65 ;
        RECT  0.50 5.00 4.45 5.50 ;
        RECT  3.75 5.00 4.45 5.70 ;
        RECT  4.20 3.55 5.40 4.25 ;
        RECT  4.20 8.65 4.90 10.25 ;
        RECT  4.90 3.55 5.40 9.15 ;
        RECT  4.20 8.65 5.40 9.15 ;
        RECT  7.75 2.55 8.25 5.10 ;
        RECT  4.90 4.60 8.25 5.10 ;
        RECT  8.90 3.55 9.60 4.25 ;
        RECT  9.10 3.55 9.60 10.00 ;
        RECT  8.90 8.40 9.60 10.00 ;
        RECT  7.75 2.55 10.70 3.05 ;
        RECT  10.20 2.55 10.70 5.10 ;
        RECT  10.20 4.60 12.40 5.10 ;
        RECT  11.70 4.60 12.40 5.30 ;
        RECT  13.60 3.55 14.30 5.25 ;
        RECT  13.60 7.40 14.30 10.05 ;
        RECT  9.10 5.75 15.40 6.25 ;
        RECT  14.70 5.75 15.40 6.45 ;
        RECT  13.60 4.75 16.40 5.25 ;
        RECT  15.90 4.75 16.40 7.90 ;
        RECT  13.60 7.40 16.40 7.90 ;
        RECT  17.30 8.30 18.00 10.05 ;
        RECT  17.70 5.55 18.40 6.25 ;
        RECT  15.90 5.75 18.40 6.25 ;
        RECT  17.30 3.55 19.35 4.25 ;
        RECT  18.85 3.55 19.35 8.80 ;
        RECT  17.30 8.30 19.35 8.80 ;
    END
END MU4IX4
MACRO MU4X1
    CLASS CORE ;
    FOREIGN MU4X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN S1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.40 19.35 6.30 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  0.25 6.70 1.25 7.60 ;
        END
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M2M ;
        RECT  14.35 2.85 15.05 9.00 ;
        RECT  14.30 2.85 15.10 3.65 ;
        RECT  14.30 7.90 15.10 9.00 ;
        LAYER M1M ;
        RECT  14.25 2.45 15.15 4.05 ;
        RECT  14.25 7.55 15.15 10.45 ;
        END
    END Q
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.20 6.70 8.15 7.60 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  10.05 6.70 10.95 7.60 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 6.70 6.75 7.60 ;
        END
    END IN1
    PIN IN0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END IN0
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 9.55 2.50 11.00 ;
        RECT  6.50 8.60 7.20 11.00 ;
        RECT  11.20 8.60 12.80 10.20 ;
        RECT  12.10 7.25 12.80 11.00 ;
        RECT  16.80 7.75 17.50 11.00 ;
        RECT  18.45 10.10 19.15 11.00 ;
        RECT  0.00 11.00 19.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.05 ;
        RECT  6.50 2.00 7.20 4.00 ;
        RECT  11.20 2.00 12.80 4.00 ;
        RECT  16.80 2.00 17.50 4.00 ;
        RECT  0.00 0.00 19.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.35 1.15 4.05 ;
        RECT  0.65 3.35 1.15 5.40 ;
        RECT  0.45 8.15 1.15 10.25 ;
        RECT  1.75 4.90 2.25 8.65 ;
        RECT  0.45 8.15 2.25 8.65 ;
        RECT  3.70 4.70 4.40 5.40 ;
        RECT  0.65 4.90 4.40 5.40 ;
        RECT  4.15 3.35 5.35 4.05 ;
        RECT  4.15 8.60 4.85 10.20 ;
        RECT  4.85 3.35 5.35 9.10 ;
        RECT  4.15 8.60 5.35 9.10 ;
        RECT  7.70 2.45 8.20 5.40 ;
        RECT  4.85 4.90 8.20 5.40 ;
        RECT  8.85 3.40 9.55 4.10 ;
        RECT  9.05 3.40 9.55 10.20 ;
        RECT  8.85 8.60 9.55 10.20 ;
        RECT  7.70 2.45 10.60 2.95 ;
        RECT  10.10 2.45 10.60 5.00 ;
        RECT  10.10 4.50 13.25 5.00 ;
        RECT  12.55 4.50 13.25 5.20 ;
        RECT  13.80 4.95 14.30 6.15 ;
        RECT  9.05 5.65 14.30 6.15 ;
        RECT  14.90 5.90 15.60 6.60 ;
        RECT  16.15 4.75 16.85 5.45 ;
        RECT  13.80 4.95 16.85 5.45 ;
        RECT  14.90 6.10 17.80 6.60 ;
        RECT  17.30 4.45 17.80 7.25 ;
        RECT  17.30 6.75 19.00 7.25 ;
        RECT  18.30 3.40 19.00 4.95 ;
        RECT  17.30 4.45 19.00 4.95 ;
        RECT  18.30 6.75 19.00 8.85 ;
        LAYER V1M ;
        RECT  14.20 7.95 15.20 8.95 ;
        RECT  14.20 2.75 15.20 3.75 ;
    END
END MU4X1
MACRO MU4X2
    CLASS CORE ;
    FOREIGN MU4X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 28.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN S1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.25 ;
        PORT
        LAYER M1M ;
        RECT  26.85 5.40 27.75 6.30 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  0.25 6.70 1.25 7.60 ;
        END
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M2M ;
        RECT  18.55 2.50 19.25 7.70 ;
        RECT  18.50 2.50 19.30 3.30 ;
        RECT  18.50 6.60 19.30 7.70 ;
        LAYER M1M ;
        RECT  15.60 2.45 16.30 3.70 ;
        RECT  15.60 7.75 16.30 10.55 ;
        RECT  18.30 2.45 19.00 4.50 ;
        RECT  18.45 6.65 19.00 10.55 ;
        RECT  18.30 7.10 19.00 10.55 ;
        RECT  18.30 2.45 19.35 3.35 ;
        RECT  18.45 6.65 19.35 7.60 ;
        RECT  18.30 7.10 19.35 7.60 ;
        RECT  15.60 2.45 21.70 2.95 ;
        RECT  21.00 2.45 21.70 3.70 ;
        RECT  21.00 8.70 21.70 10.55 ;
        RECT  15.60 10.05 21.70 10.55 ;
        END
    END Q
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.20 6.70 8.15 7.60 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  10.05 6.70 10.95 7.60 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 6.70 6.75 7.60 ;
        END
    END IN1
    PIN IN0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END IN0
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 9.55 2.50 11.00 ;
        RECT  6.50 8.60 7.20 11.00 ;
        RECT  11.40 7.25 12.10 11.00 ;
        RECT  14.10 7.75 14.80 11.00 ;
        RECT  22.50 8.65 23.20 11.00 ;
        RECT  25.20 7.70 25.90 11.00 ;
        RECT  26.85 10.25 27.55 11.00 ;
        RECT  0.00 11.00 28.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.05 ;
        RECT  6.50 2.00 7.20 4.00 ;
        RECT  11.40 2.00 12.10 4.15 ;
        RECT  14.10 2.00 14.80 3.70 ;
        RECT  22.50 2.00 23.20 3.70 ;
        RECT  25.20 2.00 25.90 3.95 ;
        RECT  0.00 0.00 28.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.35 1.15 4.05 ;
        RECT  0.65 3.35 1.15 5.40 ;
        RECT  0.45 8.15 1.15 10.25 ;
        RECT  1.75 4.90 2.25 8.65 ;
        RECT  0.45 8.15 2.25 8.65 ;
        RECT  3.70 4.70 4.40 5.40 ;
        RECT  0.65 4.90 4.40 5.40 ;
        RECT  4.15 3.35 5.35 4.05 ;
        RECT  4.15 8.60 4.85 10.20 ;
        RECT  4.85 3.35 5.35 9.10 ;
        RECT  4.15 8.60 5.35 9.10 ;
        RECT  7.70 2.45 8.20 5.40 ;
        RECT  4.85 4.90 8.20 5.40 ;
        RECT  8.85 3.40 9.55 4.10 ;
        RECT  9.05 3.40 9.55 10.20 ;
        RECT  8.85 8.60 9.55 10.20 ;
        RECT  7.70 2.45 10.60 2.95 ;
        RECT  10.10 2.45 10.60 5.10 ;
        RECT  10.10 4.60 12.30 5.10 ;
        RECT  11.60 4.60 12.30 5.30 ;
        RECT  12.80 5.10 13.30 6.25 ;
        RECT  9.05 5.75 13.30 6.25 ;
        RECT  12.75 2.45 13.45 4.65 ;
        RECT  12.75 6.80 13.45 10.55 ;
        RECT  12.75 6.80 17.65 7.30 ;
        RECT  16.95 3.45 17.65 4.65 ;
        RECT  12.75 4.15 17.65 4.65 ;
        RECT  16.95 6.80 17.65 9.60 ;
        RECT  19.65 3.70 20.35 4.65 ;
        RECT  19.80 7.70 20.35 9.60 ;
        RECT  19.65 7.95 20.35 9.60 ;
        RECT  22.10 6.05 22.80 6.75 ;
        RECT  12.80 5.10 24.10 5.60 ;
        RECT  19.80 7.70 24.55 8.20 ;
        RECT  19.65 7.95 24.55 8.20 ;
        RECT  23.40 5.10 24.10 5.80 ;
        RECT  23.85 2.70 24.55 4.65 ;
        RECT  19.65 4.15 24.55 4.65 ;
        RECT  23.85 7.70 24.55 10.55 ;
        RECT  25.70 4.45 26.20 7.25 ;
        RECT  22.10 6.25 26.20 6.75 ;
        RECT  25.70 6.75 27.40 7.25 ;
        RECT  26.70 3.40 27.40 4.95 ;
        RECT  25.70 4.45 27.40 4.95 ;
        RECT  26.70 6.75 27.40 8.85 ;
        LAYER V1M ;
        RECT  18.40 6.65 19.40 7.65 ;
        RECT  18.40 2.75 19.40 3.75 ;
    END
END MU4X2
MACRO MU4X4
    CLASS CORE ;
    FOREIGN MU4X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 39.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN S1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 10.50 ;
        PORT
        LAYER M1M ;
        RECT  38.05 5.40 38.95 6.30 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.25 ;
        PORT
        LAYER M1M ;
        RECT  1.45 5.40 2.55 6.30 ;
        END
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M2M ;
        RECT  24.15 2.50 24.85 7.70 ;
        RECT  24.10 2.50 24.90 3.30 ;
        RECT  24.10 6.60 24.90 7.70 ;
        LAYER M1M ;
        RECT  18.70 2.45 19.40 3.70 ;
        RECT  18.70 7.75 19.40 10.55 ;
        RECT  21.40 2.45 22.10 3.70 ;
        RECT  21.40 7.75 22.10 10.55 ;
        RECT  24.05 2.45 24.80 4.50 ;
        RECT  24.10 6.70 24.80 10.55 ;
        RECT  24.05 2.45 24.95 3.35 ;
        RECT  24.05 6.70 24.95 7.60 ;
        RECT  26.80 2.45 27.50 3.70 ;
        RECT  26.80 8.15 27.50 10.55 ;
        RECT  18.70 2.45 30.20 2.95 ;
        RECT  29.50 2.45 30.20 3.70 ;
        RECT  29.50 8.15 30.20 10.55 ;
        RECT  18.70 10.05 30.20 10.55 ;
        END
    END Q
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  10.90 5.40 12.35 6.30 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.80 6.30 ;
        END
    END IN1
    PIN IN0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END IN0
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.15 7.15 2.85 11.00 ;
        RECT  7.10 7.90 7.80 11.00 ;
        RECT  11.80 8.10 12.50 11.00 ;
        RECT  14.50 8.60 15.20 11.00 ;
        RECT  17.20 7.75 17.90 11.00 ;
        RECT  31.00 8.15 31.70 11.00 ;
        RECT  33.70 8.15 34.40 11.00 ;
        RECT  36.40 7.70 37.10 11.00 ;
        RECT  0.00 11.00 39.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.40 2.00 3.10 4.00 ;
        RECT  7.10 2.00 7.80 3.75 ;
        RECT  11.80 2.00 12.50 3.70 ;
        RECT  14.50 2.00 15.20 3.15 ;
        RECT  17.20 2.00 17.90 3.70 ;
        RECT  31.00 2.00 31.70 3.70 ;
        RECT  33.70 2.00 34.40 3.70 ;
        RECT  36.40 2.00 37.10 3.95 ;
        RECT  0.00 0.00 39.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.75 3.45 5.85 3.95 ;
        RECT  13.15 3.60 14.45 4.00 ;
        RECT  10.85 4.60 13.50 4.95 ;
        RECT  0.30 2.45 1.00 3.15 ;
        RECT  0.50 2.45 1.00 8.90 ;
        RECT  0.50 7.10 1.25 8.90 ;
        RECT  0.50 3.50 1.60 4.95 ;
        RECT  0.50 4.45 4.90 4.95 ;
        RECT  4.40 4.45 4.90 6.10 ;
        RECT  4.40 5.40 5.10 6.10 ;
        RECT  4.50 6.75 5.20 10.55 ;
        RECT  5.35 3.25 5.45 4.95 ;
        RECT  4.75 3.25 5.45 3.95 ;
        RECT  5.35 3.45 5.85 4.95 ;
        RECT  5.35 4.45 9.10 4.95 ;
        RECT  8.60 2.45 9.00 7.25 ;
        RECT  8.50 2.45 9.00 4.95 ;
        RECT  8.60 4.45 9.10 7.25 ;
        RECT  4.50 6.75 9.10 7.25 ;
        RECT  9.45 3.40 10.15 4.10 ;
        RECT  9.65 3.40 10.15 10.55 ;
        RECT  9.45 8.05 10.15 10.55 ;
        RECT  8.50 2.45 11.35 2.95 ;
        RECT  10.85 2.45 11.35 4.95 ;
        RECT  12.80 4.45 13.30 5.30 ;
        RECT  10.85 4.45 13.30 4.95 ;
        RECT  12.80 5.75 13.30 7.25 ;
        RECT  9.65 6.75 13.30 7.25 ;
        RECT  12.80 4.60 13.50 5.30 ;
        RECT  13.60 3.25 13.85 4.10 ;
        RECT  13.15 3.25 13.85 4.00 ;
        RECT  13.75 6.80 13.85 10.55 ;
        RECT  13.15 7.70 13.85 10.55 ;
        RECT  13.60 3.50 14.20 4.10 ;
        RECT  13.60 3.60 14.45 4.10 ;
        RECT  13.95 3.50 14.20 4.65 ;
        RECT  13.15 3.50 14.20 4.00 ;
        RECT  13.75 6.80 14.25 8.20 ;
        RECT  13.15 7.70 14.25 8.20 ;
        RECT  13.95 3.60 14.45 4.65 ;
        RECT  13.95 5.10 14.45 6.25 ;
        RECT  12.80 5.75 14.45 6.25 ;
        RECT  15.85 2.45 16.55 4.65 ;
        RECT  15.85 6.80 16.55 10.55 ;
        RECT  20.05 3.40 20.75 4.65 ;
        RECT  20.05 6.80 20.75 9.60 ;
        RECT  13.75 6.80 23.45 7.30 ;
        RECT  22.75 3.45 23.45 4.65 ;
        RECT  13.95 4.15 23.45 4.65 ;
        RECT  22.75 6.80 23.45 9.60 ;
        RECT  25.45 3.45 26.15 4.65 ;
        RECT  25.60 7.20 26.15 9.60 ;
        RECT  25.45 7.95 26.15 9.60 ;
        RECT  28.15 3.40 28.85 4.65 ;
        RECT  28.15 7.20 28.85 9.60 ;
        RECT  30.65 6.05 31.35 6.75 ;
        RECT  13.95 5.10 32.60 5.60 ;
        RECT  31.90 5.10 32.60 5.80 ;
        RECT  32.35 2.70 33.05 4.65 ;
        RECT  32.35 7.20 33.05 10.55 ;
        RECT  25.60 7.20 35.75 7.70 ;
        RECT  35.05 2.70 35.75 4.65 ;
        RECT  25.45 4.15 35.75 4.65 ;
        RECT  35.05 7.20 35.75 10.55 ;
        RECT  36.90 4.45 37.40 7.25 ;
        RECT  30.65 6.25 37.40 6.75 ;
        RECT  36.90 6.75 38.60 7.25 ;
        RECT  37.90 2.70 38.60 4.95 ;
        RECT  36.90 4.45 38.60 4.95 ;
        RECT  37.90 6.75 38.60 10.50 ;
        LAYER V1M ;
        RECT  24.00 6.65 25.00 7.65 ;
        RECT  24.00 2.75 25.00 3.75 ;
    END
END MU4X4
MACRO MU8IX1
    CLASS CORE ;
    FOREIGN MU8IX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 46.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN S2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  20.50 5.60 21.20 8.35 ;
        RECT  20.50 6.55 22.15 7.60 ;
        END
    END S2
    PIN S1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  16.85 8.00 17.95 8.90 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.25 ;
        PORT
        LAYER M1M ;
        RECT  1.45 6.70 2.55 7.60 ;
        END
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M2M ;
        RECT  28.30 2.85 29.10 10.30 ;
        LAYER M1M ;
        RECT  28.25 8.95 29.15 10.55 ;
        RECT  28.25 2.80 29.65 3.90 ;
        END
    END Q
    PIN IN7
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  39.45 6.70 40.35 7.60 ;
        END
    END IN7
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  35.25 8.00 36.20 8.90 ;
        END
    END IN6
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  40.85 6.70 41.75 7.60 ;
        END
    END IN5
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  43.65 5.40 44.60 6.30 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 6.70 8.15 7.60 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  10.95 8.00 12.35 8.90 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 6.70 6.75 7.60 ;
        END
    END IN1
    PIN IN0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END IN0
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.55 2.50 11.00 ;
        RECT  6.55 8.55 7.25 11.00 ;
        RECT  11.50 10.30 12.20 11.00 ;
        RECT  16.40 9.35 17.10 11.00 ;
        RECT  20.80 9.80 21.50 11.00 ;
        RECT  25.55 8.90 26.25 11.00 ;
        RECT  29.85 9.20 30.55 11.00 ;
        RECT  34.85 10.30 35.55 11.00 ;
        RECT  39.85 8.55 40.55 11.00 ;
        RECT  44.55 8.55 45.25 11.00 ;
        RECT  0.00 11.00 46.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  21.05 4.65 22.35 5.15 ;
        RECT  1.80 2.00 2.50 4.35 ;
        RECT  6.55 2.00 7.25 4.35 ;
        RECT  11.60 2.00 12.30 4.35 ;
        RECT  16.85 2.00 17.55 4.35 ;
        RECT  21.65 2.00 21.75 6.05 ;
        RECT  21.05 2.00 21.75 5.15 ;
        RECT  21.65 4.65 22.35 6.05 ;
        RECT  20.00 2.00 26.60 3.25 ;
        RECT  26.10 2.00 26.60 6.00 ;
        RECT  26.10 5.30 27.05 6.00 ;
        RECT  30.30 2.00 31.00 3.90 ;
        RECT  35.00 2.00 35.70 3.90 ;
        RECT  39.85 2.00 40.55 4.35 ;
        RECT  44.55 2.00 45.25 4.40 ;
        RECT  0.00 0.00 46.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.70 0.95 10.15 ;
        RECT  0.45 3.70 1.15 5.55 ;
        RECT  0.45 8.55 1.15 10.15 ;
        RECT  0.45 5.05 4.40 5.55 ;
        RECT  3.70 5.05 4.40 5.75 ;
        RECT  4.15 3.70 5.35 4.40 ;
        RECT  4.40 6.70 4.90 10.15 ;
        RECT  4.85 3.70 4.90 10.15 ;
        RECT  4.15 8.55 4.90 10.15 ;
        RECT  4.85 3.70 5.35 7.20 ;
        RECT  4.40 6.70 5.35 7.20 ;
        RECT  8.55 5.75 9.25 6.45 ;
        RECT  8.75 5.75 9.25 8.75 ;
        RECT  4.85 4.80 10.20 5.30 ;
        RECT  9.00 9.35 9.70 10.05 ;
        RECT  9.70 4.80 10.20 6.65 ;
        RECT  8.75 8.05 10.35 8.75 ;
        RECT  9.00 3.65 11.15 4.35 ;
        RECT  10.65 3.65 11.15 5.35 ;
        RECT  9.70 5.95 12.40 6.65 ;
        RECT  10.65 4.85 13.35 5.35 ;
        RECT  12.85 2.55 13.35 9.85 ;
        RECT  9.00 9.35 13.35 9.85 ;
        RECT  13.80 5.95 14.50 8.85 ;
        RECT  13.95 3.70 15.45 4.40 ;
        RECT  13.80 8.15 15.00 8.85 ;
        RECT  14.95 3.70 15.45 7.55 ;
        RECT  12.85 2.55 16.40 3.05 ;
        RECT  15.45 7.05 15.95 10.45 ;
        RECT  13.95 9.75 15.95 10.45 ;
        RECT  15.90 2.55 16.40 5.50 ;
        RECT  15.90 4.80 16.60 5.50 ;
        RECT  17.45 6.85 18.15 7.55 ;
        RECT  14.95 7.05 18.15 7.55 ;
        RECT  18.20 3.70 19.10 4.40 ;
        RECT  18.40 8.15 18.90 10.45 ;
        RECT  18.60 3.70 18.90 10.45 ;
        RECT  17.75 9.75 18.90 10.45 ;
        RECT  18.60 3.70 19.10 8.90 ;
        RECT  18.40 8.15 19.10 8.90 ;
        RECT  19.55 4.45 20.05 10.05 ;
        RECT  19.55 8.80 20.15 10.05 ;
        RECT  19.45 9.35 20.15 10.05 ;
        RECT  19.55 4.45 20.40 5.15 ;
        RECT  22.10 8.25 22.60 9.30 ;
        RECT  19.55 8.80 22.60 9.30 ;
        RECT  23.35 6.85 24.05 8.75 ;
        RECT  22.10 8.25 24.05 8.75 ;
        RECT  24.00 5.30 25.05 6.00 ;
        RECT  24.55 5.30 25.05 10.00 ;
        RECT  23.20 9.30 25.05 10.00 ;
        RECT  24.55 6.85 27.45 7.35 ;
        RECT  26.75 6.85 27.45 7.55 ;
        RECT  26.90 8.00 27.60 10.50 ;
        RECT  27.10 3.55 27.80 4.85 ;
        RECT  27.70 5.30 28.40 6.00 ;
        RECT  27.90 5.30 28.40 8.50 ;
        RECT  27.90 7.80 29.55 8.50 ;
        RECT  26.90 8.00 29.55 8.50 ;
        RECT  30.00 4.35 30.50 8.75 ;
        RECT  30.95 5.60 31.65 6.30 ;
        RECT  31.10 6.80 31.80 7.55 ;
        RECT  30.00 8.25 32.90 8.75 ;
        RECT  32.20 8.25 32.90 10.45 ;
        RECT  32.65 3.20 33.35 4.85 ;
        RECT  27.10 4.35 33.35 4.85 ;
        RECT  33.15 6.60 33.85 7.30 ;
        RECT  31.10 6.80 33.85 7.30 ;
        RECT  34.30 5.60 34.80 9.85 ;
        RECT  36.25 2.55 36.75 5.05 ;
        RECT  34.40 4.35 36.75 5.05 ;
        RECT  34.30 9.35 38.20 9.85 ;
        RECT  37.20 3.65 37.70 6.10 ;
        RECT  30.95 5.60 37.70 6.10 ;
        RECT  37.20 3.65 38.20 4.35 ;
        RECT  37.50 9.35 38.20 10.20 ;
        RECT  38.15 5.75 38.65 8.80 ;
        RECT  36.80 8.10 38.65 8.80 ;
        RECT  38.15 5.75 38.85 6.45 ;
        RECT  36.25 2.55 39.40 3.05 ;
        RECT  38.90 2.55 39.40 5.30 ;
        RECT  42.20 3.70 42.90 5.30 ;
        RECT  38.90 4.80 42.90 5.30 ;
        RECT  42.40 3.70 42.90 10.15 ;
        RECT  42.20 8.55 42.90 10.15 ;
        LAYER V1M ;
        RECT  28.20 9.25 29.20 10.25 ;
        RECT  28.20 2.75 29.20 3.75 ;
    END
END MU8IX1
MACRO MU8IX2
    CLASS CORE ;
    FOREIGN MU8IX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 46.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN S2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  20.50 5.50 21.20 8.35 ;
        RECT  20.50 6.70 22.15 7.60 ;
        END
    END S2
    PIN S1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  16.85 8.00 17.95 8.90 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.25 ;
        PORT
        LAYER M1M ;
        RECT  1.45 6.70 2.55 7.60 ;
        END
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M2M ;
        RECT  28.40 4.05 29.00 10.30 ;
        RECT  28.30 4.05 29.10 4.85 ;
        RECT  28.30 9.20 29.10 10.30 ;
        LAYER M1M ;
        RECT  28.75 3.20 29.45 4.90 ;
        RECT  28.25 4.00 29.45 4.90 ;
        RECT  28.70 7.80 29.45 10.55 ;
        RECT  28.25 9.30 29.45 10.55 ;
        END
    END Q
    PIN IN7
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  39.45 6.70 40.35 7.60 ;
        END
    END IN7
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  36.65 6.70 37.55 7.60 ;
        RECT  35.80 6.90 37.55 7.60 ;
        END
    END IN6
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  40.85 6.70 41.75 7.60 ;
        END
    END IN5
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  43.65 5.40 44.60 6.30 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 6.70 8.15 7.60 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  10.95 8.00 12.35 8.90 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 6.70 6.75 7.60 ;
        END
    END IN1
    PIN IN0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END IN0
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.55 2.50 11.00 ;
        RECT  6.55 8.55 7.25 11.00 ;
        RECT  11.50 10.30 12.20 11.00 ;
        RECT  16.40 9.35 17.10 11.00 ;
        RECT  20.80 9.80 21.50 11.00 ;
        RECT  25.55 8.90 26.25 11.00 ;
        RECT  30.10 9.20 30.80 11.00 ;
        RECT  35.00 10.30 35.70 11.00 ;
        RECT  39.85 8.55 40.55 11.00 ;
        RECT  44.55 8.55 45.25 11.00 ;
        RECT  0.00 11.00 46.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.35 ;
        RECT  6.55 2.00 7.25 4.35 ;
        RECT  11.60 2.00 12.30 4.35 ;
        RECT  16.85 2.00 17.55 4.35 ;
        RECT  21.05 2.00 21.75 5.05 ;
        RECT  25.75 2.00 26.45 5.00 ;
        RECT  30.10 2.00 30.80 4.45 ;
        RECT  35.00 2.00 35.70 3.90 ;
        RECT  39.85 2.00 40.55 4.35 ;
        RECT  44.55 2.00 45.25 4.40 ;
        RECT  0.00 0.00 46.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.70 0.95 10.15 ;
        RECT  0.45 3.70 1.15 5.55 ;
        RECT  0.45 8.55 1.15 10.15 ;
        RECT  0.45 5.05 4.40 5.55 ;
        RECT  3.70 5.05 4.40 5.75 ;
        RECT  4.15 3.70 5.35 4.40 ;
        RECT  4.40 6.70 4.90 10.15 ;
        RECT  4.85 3.70 4.90 10.15 ;
        RECT  4.15 8.55 4.90 10.15 ;
        RECT  4.85 3.70 5.35 7.20 ;
        RECT  4.40 6.70 5.35 7.20 ;
        RECT  8.55 5.75 9.25 6.45 ;
        RECT  8.75 5.75 9.25 8.75 ;
        RECT  4.85 4.80 10.20 5.30 ;
        RECT  9.00 9.35 9.70 10.05 ;
        RECT  9.70 4.80 10.20 6.65 ;
        RECT  8.75 8.05 10.35 8.75 ;
        RECT  9.00 3.65 11.15 4.35 ;
        RECT  10.65 3.65 11.15 5.35 ;
        RECT  9.70 5.95 12.40 6.65 ;
        RECT  10.65 4.85 13.35 5.35 ;
        RECT  12.85 2.55 13.35 9.85 ;
        RECT  9.00 9.35 13.35 9.85 ;
        RECT  13.80 5.95 14.50 8.85 ;
        RECT  13.95 3.70 15.45 4.40 ;
        RECT  13.80 8.15 15.00 8.85 ;
        RECT  14.95 3.70 15.45 7.55 ;
        RECT  12.85 2.55 16.40 3.05 ;
        RECT  15.45 7.05 15.95 10.45 ;
        RECT  13.95 9.75 15.95 10.45 ;
        RECT  15.90 2.55 16.40 5.50 ;
        RECT  15.90 4.80 16.60 5.50 ;
        RECT  17.45 6.85 18.15 7.55 ;
        RECT  14.95 7.05 18.15 7.55 ;
        RECT  18.20 3.70 19.10 4.40 ;
        RECT  18.40 8.15 18.90 10.45 ;
        RECT  18.60 3.70 18.90 10.45 ;
        RECT  17.75 9.75 18.90 10.45 ;
        RECT  18.60 3.70 19.10 8.90 ;
        RECT  18.40 8.15 19.10 8.90 ;
        RECT  19.55 4.35 20.05 10.05 ;
        RECT  19.55 8.80 20.15 10.05 ;
        RECT  19.45 9.35 20.15 10.05 ;
        RECT  19.55 4.35 20.40 5.05 ;
        RECT  22.10 8.25 22.60 9.30 ;
        RECT  19.55 8.80 22.60 9.30 ;
        RECT  22.75 6.85 23.45 8.75 ;
        RECT  22.10 8.25 23.45 8.75 ;
        RECT  23.40 4.30 24.40 5.00 ;
        RECT  23.90 4.30 24.40 10.00 ;
        RECT  23.20 9.30 24.40 10.00 ;
        RECT  23.90 6.85 26.85 7.35 ;
        RECT  26.15 6.85 26.85 7.55 ;
        RECT  27.10 4.30 27.80 5.00 ;
        RECT  27.30 4.30 27.60 10.50 ;
        RECT  26.90 8.00 27.60 10.50 ;
        RECT  27.30 4.30 27.80 8.50 ;
        RECT  26.90 8.00 27.80 8.50 ;
        RECT  28.25 5.35 28.95 6.05 ;
        RECT  28.95 6.60 29.65 7.30 ;
        RECT  27.30 6.80 29.65 7.30 ;
        RECT  28.25 5.55 31.15 6.05 ;
        RECT  30.65 4.90 31.15 8.75 ;
        RECT  31.60 5.85 32.30 6.55 ;
        RECT  31.60 7.10 32.30 7.80 ;
        RECT  30.65 8.25 33.20 8.75 ;
        RECT  32.50 8.25 33.20 10.45 ;
        RECT  32.65 3.20 33.35 5.40 ;
        RECT  30.65 4.90 33.35 5.40 ;
        RECT  31.60 7.10 34.35 7.60 ;
        RECT  33.65 7.10 34.35 7.80 ;
        RECT  31.60 5.85 35.35 6.35 ;
        RECT  34.85 5.70 35.35 9.85 ;
        RECT  36.25 2.55 36.75 5.05 ;
        RECT  34.45 4.35 36.75 5.05 ;
        RECT  34.85 5.70 37.70 6.20 ;
        RECT  34.85 9.35 38.20 9.85 ;
        RECT  37.20 3.65 37.70 6.20 ;
        RECT  31.60 5.85 37.70 6.20 ;
        RECT  37.20 3.65 38.20 4.35 ;
        RECT  37.50 9.35 38.20 10.20 ;
        RECT  38.15 5.75 38.65 8.85 ;
        RECT  36.80 8.15 38.65 8.85 ;
        RECT  38.15 5.75 38.85 6.45 ;
        RECT  36.25 2.55 39.40 3.05 ;
        RECT  38.90 2.55 39.40 5.30 ;
        RECT  42.20 3.70 42.90 5.30 ;
        RECT  38.90 4.80 42.90 5.30 ;
        RECT  42.40 3.70 42.90 10.15 ;
        RECT  42.20 8.55 42.90 10.15 ;
        LAYER V1M ;
        RECT  28.20 9.25 29.20 10.25 ;
        RECT  28.20 4.05 29.20 5.05 ;
    END
END MU8IX2
MACRO MU8IX4
    CLASS CORE ;
    FOREIGN MU8IX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 47.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN S2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  20.50 5.50 21.20 8.35 ;
        RECT  20.50 6.70 22.15 7.60 ;
        END
    END S2
    PIN S1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  16.85 8.00 17.95 8.90 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.25 ;
        PORT
        LAYER M1M ;
        RECT  1.45 6.70 2.55 7.60 ;
        END
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M2M ;
        RECT  29.80 4.35 30.40 9.00 ;
        RECT  29.70 7.90 30.50 9.00 ;
        RECT  29.80 4.35 30.60 5.15 ;
        LAYER M1M ;
        RECT  29.65 8.00 30.80 8.90 ;
        RECT  30.10 3.20 30.80 5.20 ;
        RECT  29.75 4.30 30.80 5.20 ;
        RECT  30.10 7.75 30.80 10.55 ;
        END
    END Q
    PIN IN7
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  40.85 6.70 41.75 7.60 ;
        END
    END IN7
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  38.05 6.70 38.95 7.60 ;
        RECT  37.20 6.90 38.95 7.60 ;
        END
    END IN6
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  42.25 6.70 43.15 7.60 ;
        END
    END IN5
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  45.05 5.40 46.00 6.30 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 6.70 8.15 7.60 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  10.95 8.00 12.35 8.90 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 6.70 6.75 7.60 ;
        END
    END IN1
    PIN IN0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END IN0
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.55 2.50 11.00 ;
        RECT  6.55 8.55 7.25 11.00 ;
        RECT  11.50 10.30 12.20 11.00 ;
        RECT  16.40 9.35 17.10 11.00 ;
        RECT  20.80 9.80 21.50 11.00 ;
        RECT  25.70 8.70 26.40 11.00 ;
        RECT  28.75 9.35 29.45 11.00 ;
        RECT  31.45 9.20 32.15 11.00 ;
        RECT  36.40 10.30 37.10 11.00 ;
        RECT  41.25 8.55 41.95 11.00 ;
        RECT  45.95 8.55 46.65 11.00 ;
        RECT  0.00 11.00 47.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.35 ;
        RECT  6.55 2.00 7.25 4.35 ;
        RECT  11.60 2.00 12.30 4.35 ;
        RECT  16.85 2.00 17.55 4.35 ;
        RECT  21.05 2.00 21.75 5.05 ;
        RECT  25.75 2.00 26.45 5.00 ;
        RECT  28.75 2.00 29.45 3.95 ;
        RECT  31.45 2.00 32.15 3.95 ;
        RECT  36.40 2.00 37.10 3.90 ;
        RECT  41.25 2.00 41.95 4.35 ;
        RECT  45.95 2.00 46.65 4.40 ;
        RECT  0.00 0.00 47.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.70 0.95 10.15 ;
        RECT  0.45 3.70 1.15 5.55 ;
        RECT  0.45 8.55 1.15 10.15 ;
        RECT  0.45 5.05 4.40 5.55 ;
        RECT  3.70 5.05 4.40 5.75 ;
        RECT  4.15 3.70 5.35 4.40 ;
        RECT  4.40 6.70 4.90 10.15 ;
        RECT  4.85 3.70 4.90 10.15 ;
        RECT  4.15 8.55 4.90 10.15 ;
        RECT  4.85 3.70 5.35 7.20 ;
        RECT  4.40 6.70 5.35 7.20 ;
        RECT  8.55 5.75 9.25 6.45 ;
        RECT  8.75 5.75 9.25 8.75 ;
        RECT  4.85 4.80 10.20 5.30 ;
        RECT  9.00 9.35 9.70 10.05 ;
        RECT  9.70 4.80 10.20 6.65 ;
        RECT  8.75 8.05 10.35 8.75 ;
        RECT  9.00 3.65 11.15 4.35 ;
        RECT  10.65 3.65 11.15 5.35 ;
        RECT  9.70 5.95 12.40 6.65 ;
        RECT  10.65 4.85 13.35 5.35 ;
        RECT  12.85 2.55 13.35 9.85 ;
        RECT  9.00 9.35 13.35 9.85 ;
        RECT  13.80 5.95 14.50 8.85 ;
        RECT  13.95 3.70 15.45 4.40 ;
        RECT  13.80 8.15 15.00 8.85 ;
        RECT  14.95 3.70 15.45 7.55 ;
        RECT  12.85 2.55 16.40 3.05 ;
        RECT  15.45 7.05 15.95 10.45 ;
        RECT  13.95 9.75 15.95 10.45 ;
        RECT  15.90 2.55 16.40 5.50 ;
        RECT  15.90 4.80 16.60 5.50 ;
        RECT  17.45 6.85 18.15 7.55 ;
        RECT  14.95 7.05 18.15 7.55 ;
        RECT  18.20 3.70 19.10 4.40 ;
        RECT  18.40 8.15 18.90 10.45 ;
        RECT  18.60 3.70 18.90 10.45 ;
        RECT  17.75 9.75 18.90 10.45 ;
        RECT  18.60 3.70 19.10 8.90 ;
        RECT  18.40 8.15 19.10 8.90 ;
        RECT  19.55 4.35 20.05 10.05 ;
        RECT  19.55 8.80 20.15 10.05 ;
        RECT  19.45 9.35 20.15 10.05 ;
        RECT  19.55 4.35 20.40 5.05 ;
        RECT  22.10 8.25 22.60 9.30 ;
        RECT  19.55 8.80 22.60 9.30 ;
        RECT  22.75 6.85 23.45 8.75 ;
        RECT  22.10 8.25 23.45 8.75 ;
        RECT  23.40 4.30 24.40 5.00 ;
        RECT  23.90 4.30 24.40 10.00 ;
        RECT  23.20 9.30 24.40 10.00 ;
        RECT  23.90 6.85 26.85 7.35 ;
        RECT  26.15 6.85 26.85 7.55 ;
        RECT  27.10 4.30 27.80 5.00 ;
        RECT  27.30 4.30 27.80 10.50 ;
        RECT  27.10 8.70 27.80 10.50 ;
        RECT  28.25 5.65 28.95 6.35 ;
        RECT  29.65 6.60 30.35 7.30 ;
        RECT  27.30 6.80 30.35 7.30 ;
        RECT  28.25 5.65 32.55 6.15 ;
        RECT  32.05 4.90 32.55 8.75 ;
        RECT  33.00 5.85 33.70 6.55 ;
        RECT  33.00 7.10 33.70 7.80 ;
        RECT  32.05 8.25 34.60 8.75 ;
        RECT  33.90 8.25 34.60 10.45 ;
        RECT  34.05 3.20 34.75 5.40 ;
        RECT  32.05 4.90 34.75 5.40 ;
        RECT  33.00 7.10 35.75 7.60 ;
        RECT  35.05 7.10 35.75 7.80 ;
        RECT  33.00 5.85 36.75 6.35 ;
        RECT  36.25 5.70 36.75 9.85 ;
        RECT  37.65 2.55 38.15 5.05 ;
        RECT  35.85 4.35 38.15 5.05 ;
        RECT  36.25 5.70 39.10 6.20 ;
        RECT  36.25 9.35 39.60 9.85 ;
        RECT  38.60 3.65 39.10 6.20 ;
        RECT  33.00 5.85 39.10 6.20 ;
        RECT  38.60 3.65 39.60 4.35 ;
        RECT  38.90 9.35 39.60 10.20 ;
        RECT  39.55 5.75 40.05 8.85 ;
        RECT  38.20 8.15 40.05 8.85 ;
        RECT  39.55 5.75 40.25 6.45 ;
        RECT  37.65 2.55 40.80 3.05 ;
        RECT  40.30 2.55 40.80 5.30 ;
        RECT  43.60 3.70 44.30 5.30 ;
        RECT  40.30 4.80 44.30 5.30 ;
        RECT  43.80 3.70 44.30 10.15 ;
        RECT  43.60 8.55 44.30 10.15 ;
        LAYER V1M ;
        RECT  29.60 7.95 30.60 8.95 ;
        RECT  29.60 4.05 30.60 5.05 ;
    END
END MU8IX4
MACRO MU8X1
    CLASS CORE ;
    FOREIGN MU8X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 44.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN S2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  20.50 5.60 21.20 8.35 ;
        RECT  20.50 6.55 22.15 7.60 ;
        END
    END S2
    PIN S1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  16.85 8.00 17.95 8.90 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.25 ;
        PORT
        LAYER M1M ;
        RECT  1.45 6.70 2.55 7.60 ;
        END
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  27.25 4.85 27.95 5.55 ;
        RECT  27.45 4.85 27.95 10.50 ;
        RECT  26.85 8.90 27.95 10.50 ;
        END
    END Q
    PIN IN7
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  38.05 6.70 38.95 7.60 ;
        END
    END IN7
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  33.85 8.00 34.80 8.90 ;
        END
    END IN6
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  39.45 6.70 40.35 7.60 ;
        END
    END IN5
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  42.25 5.40 43.20 6.30 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 6.70 8.15 7.60 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  10.95 8.00 12.35 8.90 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 6.70 6.75 7.60 ;
        END
    END IN1
    PIN IN0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END IN0
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.55 2.50 11.00 ;
        RECT  6.55 8.55 7.25 11.00 ;
        RECT  11.50 10.30 12.20 11.00 ;
        RECT  16.40 9.35 17.10 11.00 ;
        RECT  20.80 9.80 21.50 11.00 ;
        RECT  25.55 8.90 26.25 11.00 ;
        RECT  28.40 9.35 29.10 11.00 ;
        RECT  33.45 10.30 34.15 11.00 ;
        RECT  38.45 8.55 39.15 11.00 ;
        RECT  43.15 8.55 43.85 11.00 ;
        RECT  0.00 11.00 44.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.35 ;
        RECT  6.55 2.00 7.25 4.35 ;
        RECT  11.60 2.00 12.30 4.35 ;
        RECT  16.85 2.00 17.55 4.35 ;
        RECT  21.05 2.00 21.75 5.15 ;
        RECT  25.90 2.00 26.60 5.55 ;
        RECT  20.00 2.00 27.90 3.25 ;
        RECT  28.90 2.00 29.60 3.90 ;
        RECT  33.60 2.00 34.30 3.90 ;
        RECT  38.45 2.00 39.15 4.35 ;
        RECT  43.15 2.00 43.85 4.40 ;
        RECT  0.00 0.00 44.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.70 0.95 10.15 ;
        RECT  0.45 3.70 1.15 5.55 ;
        RECT  0.45 8.55 1.15 10.15 ;
        RECT  0.45 5.05 4.40 5.55 ;
        RECT  3.70 5.05 4.40 5.75 ;
        RECT  4.15 3.70 5.35 4.40 ;
        RECT  4.40 6.70 4.90 10.15 ;
        RECT  4.85 3.70 4.90 10.15 ;
        RECT  4.15 8.55 4.90 10.15 ;
        RECT  4.85 3.70 5.35 7.20 ;
        RECT  4.40 6.70 5.35 7.20 ;
        RECT  8.55 5.75 9.25 6.45 ;
        RECT  8.75 5.75 9.25 8.75 ;
        RECT  4.85 4.80 10.20 5.30 ;
        RECT  9.00 9.35 9.70 10.05 ;
        RECT  9.70 4.80 10.20 6.65 ;
        RECT  8.75 8.05 10.35 8.75 ;
        RECT  9.00 3.65 11.15 4.35 ;
        RECT  10.65 3.65 11.15 5.35 ;
        RECT  9.70 5.95 12.40 6.65 ;
        RECT  10.65 4.85 13.35 5.35 ;
        RECT  12.85 2.55 13.35 9.85 ;
        RECT  9.00 9.35 13.35 9.85 ;
        RECT  13.80 5.95 14.50 8.85 ;
        RECT  13.95 3.70 15.45 4.40 ;
        RECT  13.80 8.15 15.00 8.85 ;
        RECT  14.95 3.70 15.45 7.55 ;
        RECT  12.85 2.55 16.40 3.05 ;
        RECT  15.45 7.05 15.95 10.45 ;
        RECT  13.95 9.75 15.95 10.45 ;
        RECT  15.90 2.55 16.40 5.50 ;
        RECT  15.90 4.80 16.60 5.50 ;
        RECT  17.45 6.85 18.15 7.55 ;
        RECT  14.95 7.05 18.15 7.55 ;
        RECT  18.20 3.70 19.10 4.40 ;
        RECT  18.40 8.15 18.90 10.45 ;
        RECT  18.60 3.70 18.90 10.45 ;
        RECT  17.75 9.75 18.90 10.45 ;
        RECT  18.60 3.70 19.10 8.90 ;
        RECT  18.40 8.15 19.10 8.90 ;
        RECT  19.55 4.45 20.05 10.05 ;
        RECT  19.55 8.80 20.15 10.05 ;
        RECT  19.45 9.35 20.15 10.05 ;
        RECT  19.55 4.45 20.40 5.15 ;
        RECT  22.10 8.25 22.60 9.30 ;
        RECT  19.55 8.80 22.60 9.30 ;
        RECT  23.10 6.15 23.60 8.75 ;
        RECT  22.10 8.25 23.60 8.75 ;
        RECT  23.10 6.15 23.80 6.85 ;
        RECT  23.55 4.85 25.05 5.55 ;
        RECT  24.55 4.85 25.05 10.00 ;
        RECT  23.20 9.30 25.05 10.00 ;
        RECT  24.55 6.05 26.95 6.85 ;
        RECT  28.55 4.35 29.05 8.75 ;
        RECT  28.55 4.35 29.25 5.05 ;
        RECT  29.55 5.60 30.25 6.30 ;
        RECT  29.65 6.95 30.35 7.70 ;
        RECT  28.55 8.25 31.45 8.75 ;
        RECT  30.75 8.25 31.45 10.45 ;
        RECT  31.25 3.20 31.95 4.85 ;
        RECT  28.55 4.35 31.95 4.85 ;
        RECT  31.70 6.60 32.40 7.45 ;
        RECT  29.65 6.95 32.40 7.45 ;
        RECT  32.90 5.60 33.40 9.85 ;
        RECT  34.85 2.55 35.35 5.05 ;
        RECT  33.00 4.35 35.35 5.05 ;
        RECT  32.90 9.35 36.80 9.85 ;
        RECT  35.80 3.65 36.30 6.10 ;
        RECT  29.55 5.60 36.30 6.10 ;
        RECT  35.80 3.65 36.80 4.35 ;
        RECT  36.10 9.35 36.80 10.20 ;
        RECT  36.75 5.75 37.25 8.80 ;
        RECT  35.40 8.10 37.25 8.80 ;
        RECT  36.75 5.75 37.45 6.45 ;
        RECT  34.85 2.55 38.00 3.05 ;
        RECT  37.50 2.55 38.00 5.30 ;
        RECT  40.80 3.70 41.50 5.30 ;
        RECT  37.50 4.80 41.50 5.30 ;
        RECT  41.00 3.70 41.50 10.15 ;
        RECT  40.80 8.55 41.50 10.15 ;
    END
END MU8X1
MACRO MU8X2
    CLASS CORE ;
    FOREIGN MU8X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 44.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN S2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  20.50 5.50 21.20 8.35 ;
        RECT  20.50 6.70 22.15 7.60 ;
        END
    END S2
    PIN S1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  16.85 8.00 17.95 8.90 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.25 ;
        PORT
        LAYER M1M ;
        RECT  1.45 6.70 2.55 7.60 ;
        END
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M2M ;
        RECT  27.00 4.05 27.60 10.30 ;
        RECT  26.90 9.20 27.70 10.30 ;
        RECT  27.00 4.05 27.80 4.85 ;
        LAYER M1M ;
        RECT  27.35 3.20 28.05 4.90 ;
        RECT  26.95 4.00 28.05 4.90 ;
        RECT  27.30 7.80 28.05 10.55 ;
        RECT  26.85 9.30 28.05 10.55 ;
        END
    END Q
    PIN IN7
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  38.05 6.70 38.95 7.60 ;
        END
    END IN7
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  35.25 6.70 36.15 7.60 ;
        RECT  34.40 6.90 36.15 7.60 ;
        END
    END IN6
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  39.45 6.70 40.35 7.60 ;
        END
    END IN5
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  42.25 5.40 43.20 6.30 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 6.70 8.15 7.60 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  10.95 8.00 12.35 8.90 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 6.70 6.75 7.60 ;
        END
    END IN1
    PIN IN0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END IN0
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.55 2.50 11.00 ;
        RECT  6.55 8.55 7.25 11.00 ;
        RECT  11.50 10.30 12.20 11.00 ;
        RECT  16.40 9.35 17.10 11.00 ;
        RECT  20.80 9.80 21.50 11.00 ;
        RECT  25.55 8.90 26.25 11.00 ;
        RECT  28.70 9.20 29.40 11.00 ;
        RECT  33.60 10.30 34.30 11.00 ;
        RECT  38.45 8.55 39.15 11.00 ;
        RECT  43.15 8.55 43.85 11.00 ;
        RECT  0.00 11.00 44.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.35 ;
        RECT  6.55 2.00 7.25 4.35 ;
        RECT  11.60 2.00 12.30 4.35 ;
        RECT  16.85 2.00 17.55 4.35 ;
        RECT  21.05 2.00 21.75 5.00 ;
        RECT  25.75 2.00 26.45 4.95 ;
        RECT  28.70 2.00 29.40 4.45 ;
        RECT  33.60 2.00 34.30 3.90 ;
        RECT  38.45 2.00 39.15 4.35 ;
        RECT  43.15 2.00 43.85 4.40 ;
        RECT  0.00 0.00 44.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.70 0.95 10.15 ;
        RECT  0.45 3.70 1.15 5.55 ;
        RECT  0.45 8.55 1.15 10.15 ;
        RECT  0.45 5.05 4.40 5.55 ;
        RECT  3.70 5.05 4.40 5.75 ;
        RECT  4.15 3.70 5.35 4.40 ;
        RECT  4.40 6.70 4.90 10.15 ;
        RECT  4.85 3.70 4.90 10.15 ;
        RECT  4.15 8.55 4.90 10.15 ;
        RECT  4.85 3.70 5.35 7.20 ;
        RECT  4.40 6.70 5.35 7.20 ;
        RECT  8.55 5.75 9.25 6.45 ;
        RECT  8.75 5.75 9.25 8.75 ;
        RECT  4.85 4.80 10.20 5.30 ;
        RECT  9.00 9.35 9.70 10.05 ;
        RECT  9.70 4.80 10.20 6.65 ;
        RECT  8.75 8.05 10.35 8.75 ;
        RECT  9.00 3.65 11.15 4.35 ;
        RECT  10.65 3.65 11.15 5.35 ;
        RECT  9.70 5.95 12.40 6.65 ;
        RECT  10.65 4.85 13.35 5.35 ;
        RECT  12.85 2.55 13.35 9.85 ;
        RECT  9.00 9.35 13.35 9.85 ;
        RECT  13.80 5.95 14.50 8.85 ;
        RECT  13.95 3.70 15.45 4.40 ;
        RECT  13.80 8.15 15.00 8.85 ;
        RECT  14.95 3.70 15.45 7.55 ;
        RECT  12.85 2.55 16.40 3.05 ;
        RECT  15.45 7.05 15.95 10.45 ;
        RECT  13.95 9.75 15.95 10.45 ;
        RECT  15.90 2.55 16.40 5.50 ;
        RECT  15.90 4.80 16.60 5.50 ;
        RECT  17.45 6.85 18.15 7.55 ;
        RECT  14.95 7.05 18.15 7.55 ;
        RECT  18.20 3.70 19.10 4.40 ;
        RECT  18.40 8.15 18.90 10.45 ;
        RECT  18.60 3.70 18.90 10.45 ;
        RECT  17.75 9.75 18.90 10.45 ;
        RECT  18.60 3.70 19.10 8.90 ;
        RECT  18.40 8.15 19.10 8.90 ;
        RECT  19.55 4.30 20.05 10.05 ;
        RECT  19.55 8.80 20.15 10.05 ;
        RECT  19.45 9.35 20.15 10.05 ;
        RECT  19.55 4.30 20.40 5.00 ;
        RECT  22.10 8.25 22.60 9.30 ;
        RECT  19.55 8.80 22.60 9.30 ;
        RECT  22.75 6.85 23.45 8.75 ;
        RECT  22.10 8.25 23.45 8.75 ;
        RECT  23.40 4.25 24.40 4.95 ;
        RECT  23.90 4.25 24.40 10.00 ;
        RECT  23.20 9.30 24.40 10.00 ;
        RECT  25.10 5.40 25.80 6.10 ;
        RECT  23.90 6.60 28.30 7.10 ;
        RECT  27.55 6.60 28.30 7.30 ;
        RECT  25.10 5.60 29.75 6.10 ;
        RECT  29.25 4.90 29.75 8.75 ;
        RECT  30.20 5.85 30.90 6.55 ;
        RECT  30.20 7.10 30.90 7.80 ;
        RECT  29.25 8.25 31.80 8.75 ;
        RECT  31.10 8.25 31.80 10.45 ;
        RECT  31.25 3.20 31.95 5.40 ;
        RECT  29.25 4.90 31.95 5.40 ;
        RECT  30.20 7.10 32.95 7.60 ;
        RECT  32.25 7.10 32.95 7.80 ;
        RECT  30.20 5.85 33.95 6.35 ;
        RECT  33.45 5.70 33.95 9.85 ;
        RECT  34.85 2.55 35.35 5.05 ;
        RECT  33.05 4.35 35.35 5.05 ;
        RECT  33.45 5.70 36.30 6.20 ;
        RECT  33.45 9.35 36.80 9.85 ;
        RECT  35.80 3.65 36.30 6.20 ;
        RECT  30.20 5.85 36.30 6.20 ;
        RECT  35.80 3.65 36.80 4.35 ;
        RECT  36.10 9.35 36.80 10.20 ;
        RECT  36.75 5.75 37.25 8.85 ;
        RECT  35.40 8.15 37.25 8.85 ;
        RECT  36.75 5.75 37.45 6.45 ;
        RECT  34.85 2.55 38.00 3.05 ;
        RECT  37.50 2.55 38.00 5.30 ;
        RECT  40.80 3.70 41.50 5.30 ;
        RECT  37.50 4.80 41.50 5.30 ;
        RECT  41.00 3.70 41.50 10.15 ;
        RECT  40.80 8.55 41.50 10.15 ;
        LAYER V1M ;
        RECT  26.80 9.25 27.80 10.25 ;
        RECT  26.80 4.05 27.80 5.05 ;
    END
END MU8X2
MACRO MU8X4
    CLASS CORE ;
    FOREIGN MU8X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 44.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN S2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  20.50 5.50 21.20 8.35 ;
        RECT  20.50 6.70 22.15 7.60 ;
        END
    END S2
    PIN S1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  16.85 8.00 17.95 8.90 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.25 ;
        PORT
        LAYER M1M ;
        RECT  1.45 6.70 2.55 7.60 ;
        END
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M2M ;
        RECT  27.00 4.35 27.60 9.00 ;
        RECT  26.90 7.90 27.70 9.00 ;
        RECT  27.00 4.35 27.80 5.15 ;
        LAYER M1M ;
        RECT  26.85 8.00 28.00 8.90 ;
        RECT  27.30 3.20 28.00 5.20 ;
        RECT  26.95 4.30 28.00 5.20 ;
        RECT  27.30 7.75 28.00 10.55 ;
        END
    END Q
    PIN IN7
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  38.05 6.70 38.95 7.60 ;
        END
    END IN7
    PIN IN6
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  35.25 6.70 36.15 7.60 ;
        RECT  34.40 6.90 36.15 7.60 ;
        END
    END IN6
    PIN IN5
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  39.45 6.70 40.35 7.60 ;
        END
    END IN5
    PIN IN4
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  42.25 5.40 43.20 6.30 ;
        END
    END IN4
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 6.70 8.15 7.60 ;
        END
    END IN3
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  10.95 8.00 12.35 8.90 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 6.70 6.75 7.60 ;
        END
    END IN1
    PIN IN0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END IN0
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.55 2.50 11.00 ;
        RECT  6.55 8.55 7.25 11.00 ;
        RECT  11.50 10.30 12.20 11.00 ;
        RECT  16.40 9.35 17.10 11.00 ;
        RECT  20.80 9.80 21.50 11.00 ;
        RECT  25.70 7.75 26.40 11.00 ;
        RECT  25.70 10.70 26.55 11.00 ;
        RECT  28.65 9.20 29.35 11.00 ;
        RECT  33.60 10.30 34.30 11.00 ;
        RECT  38.45 8.55 39.15 11.00 ;
        RECT  43.15 8.55 43.85 11.00 ;
        RECT  0.00 11.00 44.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.35 ;
        RECT  6.55 2.00 7.25 4.35 ;
        RECT  11.60 2.00 12.30 4.35 ;
        RECT  16.85 2.00 17.55 4.35 ;
        RECT  21.05 2.00 21.75 5.00 ;
        RECT  25.75 2.00 26.45 5.00 ;
        RECT  25.75 2.00 26.65 3.90 ;
        RECT  28.65 2.00 29.35 3.95 ;
        RECT  33.60 2.00 34.30 3.90 ;
        RECT  38.45 2.00 39.15 4.35 ;
        RECT  43.15 2.00 43.85 4.40 ;
        RECT  0.00 0.00 44.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.70 0.95 10.15 ;
        RECT  0.45 3.70 1.15 5.55 ;
        RECT  0.45 8.55 1.15 10.15 ;
        RECT  0.45 5.05 4.40 5.55 ;
        RECT  3.70 5.05 4.40 5.75 ;
        RECT  4.15 3.70 5.35 4.40 ;
        RECT  4.40 6.70 4.90 10.15 ;
        RECT  4.85 3.70 4.90 10.15 ;
        RECT  4.15 8.55 4.90 10.15 ;
        RECT  4.85 3.70 5.35 7.20 ;
        RECT  4.40 6.70 5.35 7.20 ;
        RECT  8.55 5.75 9.25 6.45 ;
        RECT  8.75 5.75 9.25 8.75 ;
        RECT  4.85 4.80 10.20 5.30 ;
        RECT  9.00 9.35 9.70 10.05 ;
        RECT  9.70 4.80 10.20 6.65 ;
        RECT  8.75 8.05 10.35 8.75 ;
        RECT  9.00 3.65 11.15 4.35 ;
        RECT  10.65 3.65 11.15 5.35 ;
        RECT  9.70 5.95 12.40 6.65 ;
        RECT  10.65 4.85 13.35 5.35 ;
        RECT  12.85 2.55 13.35 9.85 ;
        RECT  9.00 9.35 13.35 9.85 ;
        RECT  13.80 5.95 14.50 8.85 ;
        RECT  13.95 3.70 15.45 4.40 ;
        RECT  13.80 8.15 15.00 8.85 ;
        RECT  14.95 3.70 15.45 7.55 ;
        RECT  12.85 2.55 16.40 3.05 ;
        RECT  15.45 7.05 15.95 10.45 ;
        RECT  13.95 9.75 15.95 10.45 ;
        RECT  15.90 2.55 16.40 5.50 ;
        RECT  15.90 4.80 16.60 5.50 ;
        RECT  17.45 6.85 18.15 7.55 ;
        RECT  14.95 7.05 18.15 7.55 ;
        RECT  18.20 3.70 19.10 4.40 ;
        RECT  18.40 8.15 18.90 10.45 ;
        RECT  18.60 3.70 18.90 10.45 ;
        RECT  17.75 9.75 18.90 10.45 ;
        RECT  18.60 3.70 19.10 8.90 ;
        RECT  18.40 8.15 19.10 8.90 ;
        RECT  19.55 4.30 20.05 10.05 ;
        RECT  19.55 8.80 20.15 10.05 ;
        RECT  19.45 9.35 20.15 10.05 ;
        RECT  19.55 4.30 20.40 5.00 ;
        RECT  22.10 8.25 22.60 9.30 ;
        RECT  19.55 8.80 22.60 9.30 ;
        RECT  22.75 6.85 23.45 8.75 ;
        RECT  22.10 8.25 23.45 8.75 ;
        RECT  23.40 4.25 24.40 4.95 ;
        RECT  23.90 4.25 24.40 10.00 ;
        RECT  23.20 9.30 24.40 10.00 ;
        RECT  25.10 5.65 25.80 6.35 ;
        RECT  26.85 6.60 27.55 7.30 ;
        RECT  23.90 6.80 27.55 7.30 ;
        RECT  25.10 5.65 29.75 6.15 ;
        RECT  29.25 4.90 29.75 8.75 ;
        RECT  30.20 5.85 30.90 6.55 ;
        RECT  30.20 7.10 30.90 7.80 ;
        RECT  29.25 8.25 31.80 8.75 ;
        RECT  31.10 8.25 31.80 10.45 ;
        RECT  31.25 3.20 31.95 5.40 ;
        RECT  29.25 4.90 31.95 5.40 ;
        RECT  30.20 7.10 32.95 7.60 ;
        RECT  32.25 7.10 32.95 7.80 ;
        RECT  30.20 5.85 33.95 6.35 ;
        RECT  33.45 5.70 33.95 9.85 ;
        RECT  34.85 2.55 35.35 5.05 ;
        RECT  33.05 4.35 35.35 5.05 ;
        RECT  33.45 5.70 36.30 6.20 ;
        RECT  33.45 9.35 36.80 9.85 ;
        RECT  35.80 3.65 36.30 6.20 ;
        RECT  30.20 5.85 36.30 6.20 ;
        RECT  35.80 3.65 36.80 4.35 ;
        RECT  36.10 9.35 36.80 10.20 ;
        RECT  36.75 5.75 37.25 8.85 ;
        RECT  35.40 8.15 37.25 8.85 ;
        RECT  36.75 5.75 37.45 6.45 ;
        RECT  34.85 2.55 38.00 3.05 ;
        RECT  37.50 2.55 38.00 5.30 ;
        RECT  40.80 3.70 41.50 5.30 ;
        RECT  37.50 4.80 41.50 5.30 ;
        RECT  41.00 3.70 41.50 10.15 ;
        RECT  40.80 8.55 41.50 10.15 ;
        LAYER V1M ;
        RECT  26.80 7.95 27.80 8.95 ;
        RECT  26.80 4.05 27.80 5.05 ;
    END
END MU8X4
MACRO NA2I1X1
    CLASS CORE ;
    FOREIGN NA2I1X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.45 1.15 6.30 ;
        RECT  0.25 5.40 1.15 6.30 ;
        RECT  0.65 2.45 1.15 8.65 ;
        RECT  0.65 8.15 2.50 8.65 ;
        RECT  1.80 8.15 2.50 10.10 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.85 7.65 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 9.10 1.15 11.00 ;
        RECT  3.30 9.65 4.00 11.00 ;
        RECT  0.00 11.00 5.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.90 2.00 3.60 4.00 ;
        RECT  0.00 0.00 5.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.60 5.55 2.30 6.25 ;
        RECT  1.60 5.55 4.00 6.05 ;
        RECT  3.50 4.45 4.00 7.25 ;
        RECT  3.50 6.75 5.15 7.25 ;
        RECT  4.45 3.45 5.15 4.95 ;
        RECT  3.50 4.45 5.15 4.95 ;
        RECT  4.45 6.75 5.15 9.00 ;
    END
END NA2I1X1
MACRO NA2I1X2
    CLASS CORE ;
    FOREIGN NA2I1X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.25 6.70 1.15 7.60 ;
        RECT  0.65 2.85 0.90 8.65 ;
        RECT  0.40 2.85 0.90 7.60 ;
        RECT  0.40 2.85 1.15 4.50 ;
        RECT  0.65 6.70 1.15 8.65 ;
        RECT  0.65 8.15 2.50 8.65 ;
        RECT  1.80 8.15 2.50 10.55 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.80 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.85 7.65 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 9.10 1.15 11.00 ;
        RECT  3.15 9.50 3.85 11.00 ;
        RECT  0.00 11.00 5.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.95 2.00 3.65 4.00 ;
        RECT  0.00 0.00 5.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.35 5.55 2.05 6.25 ;
        RECT  1.35 5.55 4.00 6.05 ;
        RECT  3.50 4.45 4.00 7.25 ;
        RECT  3.50 6.75 5.15 7.25 ;
        RECT  4.45 3.75 5.15 4.95 ;
        RECT  3.50 4.45 5.15 4.95 ;
        RECT  4.45 6.75 5.15 8.85 ;
    END
END NA2I1X2
MACRO NA2I1X4
    CLASS CORE ;
    FOREIGN NA2I1X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.45 1.15 3.90 ;
        RECT  3.05 3.20 3.55 10.55 ;
        RECT  3.05 6.80 3.80 10.55 ;
        RECT  3.05 6.80 3.95 8.90 ;
        RECT  0.45 3.20 5.65 3.90 ;
        RECT  3.05 6.80 6.50 7.30 ;
        RECT  5.80 6.80 6.50 10.55 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.60 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.35 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.45 6.35 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.75 7.30 2.45 11.00 ;
        RECT  4.45 7.75 5.15 11.00 ;
        RECT  7.15 7.30 7.85 11.00 ;
        RECT  8.65 10.05 9.35 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  7.30 2.00 8.00 4.00 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.00 4.45 4.70 5.55 ;
        RECT  8.65 3.35 9.40 4.95 ;
        RECT  4.00 4.45 9.40 4.95 ;
        RECT  8.90 3.35 9.40 8.95 ;
        RECT  8.65 7.30 9.40 8.95 ;
    END
END NA2I1X4
MACRO NA2X1
    CLASS CORE ;
    FOREIGN NA2X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.65 2.75 1.35 4.60 ;
        RECT  0.65 4.10 2.55 4.60 ;
        RECT  1.60 4.10 2.10 9.15 ;
        RECT  1.60 4.10 2.55 5.00 ;
        RECT  1.60 8.45 2.65 9.15 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.50 0.75 10.20 ;
        RECT  0.25 5.50 1.05 6.20 ;
        RECT  0.25 9.30 1.15 10.20 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.55 7.10 3.60 7.80 ;
        RECT  3.10 7.10 3.60 11.00 ;
        RECT  1.60 9.80 3.60 11.00 ;
        RECT  0.00 11.00 4.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.00 2.00 3.70 4.45 ;
        RECT  0.00 0.00 4.20 2.00 ;
        END
    END gnd!
END NA2X1
MACRO NA2X2
    CLASS CORE ;
    FOREIGN NA2X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.60 2.85 1.30 4.45 ;
        RECT  0.60 3.95 2.30 4.45 ;
        RECT  1.65 8.00 2.55 8.90 ;
        RECT  1.80 3.95 2.30 10.55 ;
        RECT  1.80 7.15 2.55 10.55 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.80 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.80 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.15 1.15 11.00 ;
        RECT  3.15 7.15 3.85 11.00 ;
        RECT  0.00 11.00 5.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.95 2.00 3.65 4.40 ;
        RECT  4.45 2.00 5.15 4.70 ;
        RECT  0.00 0.00 5.60 2.00 ;
        END
    END gnd!
END NA2X2
MACRO NA2X3
    CLASS CORE ;
    FOREIGN NA2X3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.65 8.00 2.55 8.90 ;
        RECT  1.80 6.85 2.55 9.85 ;
        RECT  1.35 2.85 4.10 3.55 ;
        RECT  3.40 2.85 4.10 4.45 ;
        RECT  3.40 3.95 4.90 4.45 ;
        RECT  1.80 6.85 5.20 7.35 ;
        RECT  4.50 3.95 4.90 9.85 ;
        RECT  4.40 3.95 4.90 7.35 ;
        RECT  4.50 6.85 5.20 9.85 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.20 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.20 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.35 1.15 11.00 ;
        RECT  3.15 7.80 3.85 11.00 ;
        RECT  5.85 7.35 6.55 11.00 ;
        RECT  0.00 11.00 7.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.25 2.00 0.90 5.05 ;
        RECT  0.25 4.35 2.55 5.05 ;
        RECT  5.85 2.00 6.55 4.40 ;
        RECT  0.00 0.00 7.00 2.00 ;
        END
    END gnd!
END NA2X3
MACRO NA2X4
    CLASS CORE ;
    FOREIGN NA2X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.55 2.45 1.25 5.05 ;
        RECT  1.65 4.55 2.55 6.30 ;
        RECT  1.90 4.55 2.55 10.25 ;
        RECT  1.90 6.80 2.60 10.25 ;
        RECT  3.25 3.40 3.95 5.05 ;
        RECT  0.55 4.55 3.95 5.05 ;
        RECT  4.60 6.80 5.30 10.25 ;
        RECT  1.90 6.80 8.00 7.30 ;
        RECT  7.30 6.80 8.00 10.25 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.67 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.40 9.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.67 ;
        PORT
        LAYER M1M ;
        RECT  4.40 5.40 5.35 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.55 7.75 1.25 11.00 ;
        RECT  3.25 7.75 3.95 11.00 ;
        RECT  5.95 7.75 6.65 11.00 ;
        RECT  8.65 7.75 9.35 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  5.95 2.00 6.65 4.00 ;
        RECT  8.65 2.00 9.35 4.50 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.90 2.45 2.60 4.10 ;
        RECT  1.90 2.45 5.30 2.95 ;
        RECT  4.60 2.45 5.30 4.95 ;
        RECT  7.30 2.45 8.00 4.95 ;
        RECT  4.60 4.45 8.00 4.95 ;
    END
END NA2X4
MACRO NA3I1X1
    CLASS CORE ;
    FOREIGN NA3I1X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        RECT  1.00 2.45 1.15 9.60 ;
        RECT  0.65 4.15 1.15 9.60 ;
        RECT  0.65 7.10 1.20 9.60 ;
        RECT  0.45 7.95 1.20 9.60 ;
        RECT  1.00 2.45 1.70 4.65 ;
        RECT  0.65 4.15 1.70 4.65 ;
        RECT  0.65 7.10 3.65 7.60 ;
        RECT  3.15 7.10 3.65 9.60 ;
        RECT  3.15 7.95 3.85 9.60 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.35 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.35 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.05 2.50 11.00 ;
        RECT  4.50 8.05 5.20 11.00 ;
        RECT  0.00 11.00 7.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  4.35 2.00 5.05 4.00 ;
        RECT  0.00 0.00 7.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.15 6.90 4.85 7.60 ;
        RECT  4.90 4.45 5.40 7.40 ;
        RECT  4.15 6.90 6.35 7.40 ;
        RECT  5.85 3.80 6.35 4.95 ;
        RECT  4.90 4.45 6.35 4.95 ;
        RECT  5.85 6.90 6.35 9.60 ;
        RECT  5.85 3.80 6.55 4.50 ;
        RECT  4.90 4.45 6.55 4.50 ;
        RECT  5.85 7.95 6.55 9.60 ;
    END
END NA3I1X1
MACRO NA3I1X2
    CLASS CORE ;
    FOREIGN NA3I1X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.30 2.45 2.00 4.55 ;
        RECT  3.05 3.85 3.95 6.30 ;
        RECT  3.10 3.85 3.80 10.55 ;
        RECT  3.10 3.85 3.95 7.60 ;
        RECT  1.30 3.85 4.45 4.55 ;
        RECT  3.10 7.10 6.30 7.60 ;
        RECT  5.80 7.10 6.30 10.55 ;
        RECT  5.80 7.95 6.50 10.55 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.50 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.35 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.50 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.35 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.40 9.55 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 9.55 2.30 11.00 ;
        RECT  4.45 8.05 5.15 11.00 ;
        RECT  7.15 8.05 7.85 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  7.15 2.00 7.85 4.00 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  6.80 6.90 7.50 7.60 ;
        RECT  7.70 4.45 8.20 7.40 ;
        RECT  6.80 6.90 9.15 7.40 ;
        RECT  8.65 3.80 9.15 4.95 ;
        RECT  7.70 4.45 9.15 4.95 ;
        RECT  8.65 6.90 9.15 9.60 ;
        RECT  8.65 3.80 9.35 4.50 ;
        RECT  7.70 4.45 9.35 4.50 ;
        RECT  8.65 7.95 9.35 9.60 ;
    END
END NA3I1X2
MACRO NA3I1X4
    CLASS CORE ;
    FOREIGN NA3I1X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.90 2.45 1.60 4.80 ;
        RECT  5.85 5.40 6.75 6.30 ;
        RECT  6.25 4.10 6.70 10.55 ;
        RECT  6.00 7.10 6.70 10.55 ;
        RECT  6.25 4.10 6.75 7.60 ;
        RECT  8.70 7.10 9.40 10.55 ;
        RECT  0.90 4.10 9.95 4.80 ;
        RECT  6.00 7.10 12.10 7.60 ;
        RECT  11.40 7.10 12.10 10.55 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 7.00 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.35 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 7.00 ;
        PORT
        LAYER M1M ;
        RECT  11.30 5.40 12.35 6.35 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 9.55 3.85 11.00 ;
        RECT  4.65 8.05 5.35 11.00 ;
        RECT  7.35 8.05 8.05 11.00 ;
        RECT  10.05 8.05 10.75 11.00 ;
        RECT  12.75 8.05 13.45 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  12.75 2.00 13.45 4.00 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  13.30 4.45 13.80 7.60 ;
        RECT  12.55 6.90 13.80 7.60 ;
        RECT  12.55 7.10 14.95 7.60 ;
        RECT  14.25 3.80 14.95 4.95 ;
        RECT  13.30 4.45 14.95 4.95 ;
        RECT  14.25 7.10 14.95 9.60 ;
    END
END NA3I1X4
MACRO NA3I2X1
    CLASS CORE ;
    FOREIGN NA3I2X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        RECT  3.80 2.45 3.95 9.60 ;
        RECT  3.45 4.15 3.95 9.60 ;
        RECT  3.45 7.10 4.00 9.60 ;
        RECT  3.25 7.95 4.00 9.60 ;
        RECT  3.80 2.45 4.50 4.65 ;
        RECT  3.45 4.15 4.50 4.65 ;
        RECT  3.45 7.10 6.45 7.60 ;
        RECT  5.95 7.10 6.45 9.60 ;
        RECT  5.95 7.95 6.65 9.60 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.35 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.35 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.40 9.55 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 9.30 1.15 11.00 ;
        RECT  4.60 8.05 5.30 11.00 ;
        RECT  7.30 8.05 8.00 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 4.50 ;
        RECT  7.15 2.00 7.85 4.00 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 3.80 2.30 8.65 ;
        RECT  1.60 7.95 2.30 8.65 ;
        RECT  1.80 3.80 2.50 4.50 ;
        RECT  1.80 6.90 2.65 7.60 ;
        RECT  6.95 6.90 7.65 7.60 ;
        RECT  7.70 4.45 8.20 7.40 ;
        RECT  6.95 6.90 9.15 7.40 ;
        RECT  8.65 3.80 9.15 4.95 ;
        RECT  7.70 4.45 9.15 4.95 ;
        RECT  8.65 6.90 9.15 9.60 ;
        RECT  8.65 3.80 9.35 4.50 ;
        RECT  7.70 4.45 9.35 4.50 ;
        RECT  8.65 7.95 9.35 9.60 ;
    END
END NA3I2X1
MACRO NA3I2X2
    CLASS CORE ;
    FOREIGN NA3I2X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  2.70 2.45 3.40 4.55 ;
        RECT  4.45 3.85 5.05 10.55 ;
        RECT  4.35 6.80 5.05 10.55 ;
        RECT  4.45 3.85 5.35 7.30 ;
        RECT  2.70 3.85 5.85 4.55 ;
        RECT  4.35 6.80 7.70 7.30 ;
        RECT  7.20 6.80 7.70 10.55 ;
        RECT  7.20 7.95 7.90 10.55 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.50 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.35 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.55 7.60 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.35 8.05 2.10 11.00 ;
        RECT  5.70 7.75 6.40 11.00 ;
        RECT  8.55 8.05 9.25 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.05 2.00 1.75 3.15 ;
        RECT  8.55 2.00 9.25 4.00 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.00 3.80 1.75 4.50 ;
        RECT  1.25 3.80 1.75 5.50 ;
        RECT  1.25 5.00 3.50 5.50 ;
        RECT  3.00 5.00 3.50 9.75 ;
        RECT  2.70 8.05 3.50 9.75 ;
        RECT  3.00 6.90 3.90 7.60 ;
        RECT  8.20 6.90 8.90 7.60 ;
        RECT  9.10 4.45 9.60 7.40 ;
        RECT  8.20 6.90 10.55 7.40 ;
        RECT  10.05 3.80 10.55 4.95 ;
        RECT  9.10 4.45 10.55 4.95 ;
        RECT  10.05 6.90 10.55 9.60 ;
        RECT  10.05 3.80 10.75 4.50 ;
        RECT  9.10 4.45 10.75 4.50 ;
        RECT  10.05 7.95 10.75 9.60 ;
    END
END NA3I2X2
MACRO NA3I2X4
    CLASS CORE ;
    FOREIGN NA3I2X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  2.50 2.45 3.20 4.80 ;
        RECT  7.25 5.40 8.15 6.30 ;
        RECT  7.65 4.10 8.15 10.55 ;
        RECT  7.40 7.95 8.15 10.55 ;
        RECT  10.10 7.10 10.80 10.55 ;
        RECT  2.50 4.10 11.35 4.80 ;
        RECT  7.65 7.10 13.50 7.60 ;
        RECT  12.80 7.10 13.50 10.55 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 7.00 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.40 9.55 6.35 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.35 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 9.55 3.75 11.00 ;
        RECT  6.05 7.70 6.75 11.00 ;
        RECT  8.75 8.05 9.45 11.00 ;
        RECT  11.45 8.05 12.15 11.00 ;
        RECT  14.15 7.70 14.85 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.80 2.00 1.50 3.10 ;
        RECT  14.15 2.00 14.85 4.00 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.80 3.75 1.50 4.45 ;
        RECT  0.95 3.75 1.50 7.30 ;
        RECT  0.95 6.80 5.25 7.30 ;
        RECT  4.55 6.80 5.05 10.55 ;
        RECT  4.20 9.85 5.05 10.55 ;
        RECT  4.55 6.80 5.25 9.40 ;
        RECT  14.70 4.45 15.20 7.25 ;
        RECT  13.95 6.55 15.20 7.25 ;
        RECT  13.95 6.75 16.35 7.25 ;
        RECT  15.65 3.80 16.35 4.95 ;
        RECT  14.70 4.45 16.35 4.95 ;
        RECT  15.65 6.75 16.35 9.35 ;
    END
END NA3I2X4
MACRO NA3X1
    CLASS CORE ;
    FOREIGN NA3X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.25 2.80 1.70 3.70 ;
        RECT  0.70 2.80 1.20 10.55 ;
        RECT  1.00 2.45 1.20 10.55 ;
        RECT  0.45 8.90 1.20 10.55 ;
        RECT  1.00 2.45 1.70 4.45 ;
        RECT  0.70 2.80 1.70 4.45 ;
        RECT  0.70 8.05 3.65 8.55 ;
        RECT  3.15 8.05 3.65 10.55 ;
        RECT  3.15 8.90 3.85 10.55 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 9.00 2.50 11.00 ;
        RECT  4.50 8.95 5.20 11.00 ;
        RECT  0.00 11.00 7.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  4.35 2.00 5.05 4.50 ;
        RECT  5.85 2.00 6.55 4.70 ;
        RECT  0.00 0.00 7.00 2.00 ;
        END
    END gnd!
END NA3X1
MACRO NA3X2
    CLASS CORE ;
    FOREIGN NA3X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  2.00 5.40 2.50 10.35 ;
        RECT  1.80 9.65 2.50 10.35 ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  2.85 2.45 3.55 6.25 ;
        RECT  1.65 5.40 3.55 6.25 ;
        RECT  4.50 8.10 5.00 10.35 ;
        RECT  4.50 9.65 5.20 10.35 ;
        RECT  2.00 8.10 7.70 8.60 ;
        RECT  7.20 8.10 7.70 10.35 ;
        RECT  7.20 9.65 7.90 10.35 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.41 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.41 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.35 7.60 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.41 ;
        PORT
        LAYER M1M ;
        RECT  5.85 6.70 6.75 7.60 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 9.15 1.15 11.00 ;
        RECT  3.15 9.15 3.85 11.00 ;
        RECT  5.85 9.15 6.55 11.00 ;
        RECT  8.55 9.15 9.25 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 2.05 4.70 ;
        RECT  6.25 2.00 6.95 6.25 ;
        RECT  7.75 2.00 9.35 4.70 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
END NA3X2
MACRO NA3X3
    CLASS CORE ;
    FOREIGN NA3X3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.45 1.15 4.60 ;
        RECT  0.45 4.10 5.00 4.60 ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  2.05 4.10 2.55 8.80 ;
        RECT  3.30 8.30 4.00 10.55 ;
        RECT  2.05 4.10 5.00 4.80 ;
        RECT  4.30 4.10 5.00 6.15 ;
        RECT  6.00 8.30 6.70 10.55 ;
        RECT  2.05 8.30 9.40 8.80 ;
        RECT  8.70 8.30 9.40 10.55 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.25 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.35 7.60 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.25 ;
        PORT
        LAYER M1M ;
        RECT  5.85 6.70 6.75 7.80 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.25 ;
        PORT
        LAYER M1M ;
        RECT  8.65 6.70 9.55 7.60 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 9.55 1.15 11.00 ;
        RECT  1.95 9.25 2.65 11.00 ;
        RECT  4.65 9.25 5.35 11.00 ;
        RECT  7.35 9.25 8.05 11.00 ;
        RECT  10.05 9.25 10.75 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  7.65 2.00 8.35 6.15 ;
        RECT  9.15 2.00 10.75 4.70 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
END NA3X3
MACRO NA3X4
    CLASS CORE ;
    FOREIGN NA3X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.45 1.15 4.60 ;
        RECT  0.45 4.10 8.20 4.60 ;
        RECT  1.95 8.05 2.65 10.55 ;
        RECT  4.45 4.10 5.35 5.00 ;
        RECT  4.85 4.10 5.35 10.55 ;
        RECT  4.65 8.05 5.35 10.55 ;
        RECT  2.40 4.10 8.20 4.80 ;
        RECT  7.35 8.05 8.05 10.55 ;
        RECT  7.50 4.10 8.20 5.25 ;
        RECT  10.05 8.05 10.75 10.55 ;
        RECT  1.95 8.05 13.45 8.55 ;
        RECT  12.75 8.05 13.45 10.55 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.82 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.82 ;
        PORT
        LAYER M1M ;
        RECT  7.25 6.70 8.15 7.60 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.82 ;
        PORT
        LAYER M1M ;
        RECT  11.45 6.70 12.35 7.60 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.60 9.00 1.30 11.00 ;
        RECT  3.30 9.00 4.00 11.00 ;
        RECT  6.00 9.00 6.70 11.00 ;
        RECT  8.70 9.00 9.40 11.00 ;
        RECT  11.40 9.00 12.10 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  10.85 2.00 11.55 4.80 ;
        RECT  12.60 2.00 13.30 4.70 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
END NA3X4
MACRO NA4I1X1
    CLASS CORE ;
    FOREIGN NA4I1X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.20 3.75 10.90 4.45 ;
        RECT  10.40 3.75 10.90 8.90 ;
        RECT  10.05 7.15 10.95 8.90 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.65 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  0.25 6.70 1.15 7.60 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.25 6.50 3.95 7.60 ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 9.25 1.15 11.00 ;
        RECT  3.15 9.30 3.85 11.00 ;
        RECT  6.10 7.10 6.80 11.00 ;
        RECT  11.40 7.15 12.15 11.00 ;
        RECT  14.25 7.15 14.95 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 2.00 3.50 3.95 ;
        RECT  6.00 2.00 6.70 4.40 ;
        RECT  8.70 2.00 9.40 4.40 ;
        RECT  11.55 2.00 12.25 4.40 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.35 1.15 4.05 ;
        RECT  0.65 3.35 1.15 6.05 ;
        RECT  1.80 5.55 2.30 9.95 ;
        RECT  1.80 9.25 2.50 9.95 ;
        RECT  2.35 4.40 3.05 5.10 ;
        RECT  4.15 3.35 4.65 4.90 ;
        RECT  2.35 4.40 4.65 4.90 ;
        RECT  4.15 3.35 4.85 4.05 ;
        RECT  4.60 7.10 5.30 8.75 ;
        RECT  2.75 8.05 5.30 8.75 ;
        RECT  6.40 5.35 7.10 6.05 ;
        RECT  0.65 5.55 7.10 6.05 ;
        RECT  7.35 3.75 8.05 4.45 ;
        RECT  7.55 3.75 8.05 5.45 ;
        RECT  7.55 4.95 9.95 5.45 ;
        RECT  8.65 4.95 9.15 10.55 ;
        RECT  8.45 7.10 9.15 10.55 ;
        RECT  8.65 4.95 9.95 5.65 ;
        RECT  12.90 7.15 13.60 7.85 ;
        RECT  13.10 3.95 13.60 10.15 ;
        RECT  12.90 9.45 13.60 10.15 ;
        RECT  13.90 3.75 14.60 4.45 ;
        RECT  13.10 3.95 14.60 4.45 ;
    END
END NA4I1X1
MACRO NA4I1X2
    CLASS CORE ;
    FOREIGN NA4I1X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.20 2.70 10.90 4.50 ;
        RECT  10.40 2.70 10.90 10.55 ;
        RECT  10.05 7.10 10.95 10.55 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.70 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  0.25 6.70 1.15 7.60 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.25 6.50 3.95 7.60 ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 9.25 1.15 11.00 ;
        RECT  3.15 9.30 3.85 11.00 ;
        RECT  6.10 7.10 6.80 11.00 ;
        RECT  11.40 7.10 12.15 11.00 ;
        RECT  14.25 7.15 14.95 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 2.00 3.50 3.95 ;
        RECT  6.00 2.00 6.70 4.40 ;
        RECT  8.70 2.00 9.40 4.40 ;
        RECT  11.55 2.00 12.25 4.50 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.35 1.15 4.05 ;
        RECT  0.65 3.35 1.15 6.05 ;
        RECT  1.80 5.55 2.30 9.95 ;
        RECT  1.80 9.25 2.50 9.95 ;
        RECT  2.35 4.40 3.05 5.10 ;
        RECT  4.15 3.35 4.65 4.90 ;
        RECT  2.35 4.40 4.65 4.90 ;
        RECT  4.15 3.35 4.85 4.05 ;
        RECT  4.60 7.10 5.30 8.75 ;
        RECT  2.75 8.05 5.30 8.75 ;
        RECT  6.40 5.35 7.10 6.05 ;
        RECT  0.65 5.55 7.10 6.05 ;
        RECT  7.35 3.75 8.05 4.45 ;
        RECT  7.55 3.75 8.05 5.45 ;
        RECT  7.55 4.95 9.95 5.45 ;
        RECT  8.65 4.95 9.15 10.55 ;
        RECT  8.45 7.10 9.15 10.55 ;
        RECT  8.65 4.95 9.95 5.65 ;
        RECT  12.90 7.15 13.40 10.55 ;
        RECT  13.15 3.95 13.40 10.55 ;
        RECT  12.60 9.85 13.40 10.55 ;
        RECT  13.15 3.95 13.65 7.85 ;
        RECT  12.90 7.15 13.65 7.85 ;
        RECT  14.10 3.75 14.80 4.45 ;
        RECT  13.15 3.95 14.80 4.45 ;
    END
END NA4I1X2
MACRO NA4I1X4
    CLASS CORE ;
    FOREIGN NA4I1X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.60 2.70 12.10 10.55 ;
        RECT  11.45 7.10 12.15 10.55 ;
        RECT  11.60 2.70 12.30 4.50 ;
        RECT  11.45 7.10 12.35 8.90 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 14.10 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  0.25 6.70 1.15 7.60 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.25 6.50 3.95 7.60 ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 9.25 1.15 11.00 ;
        RECT  3.15 9.30 3.85 11.00 ;
        RECT  6.10 7.10 6.80 11.00 ;
        RECT  10.10 7.10 10.80 11.00 ;
        RECT  12.80 7.10 13.50 11.00 ;
        RECT  15.65 7.15 16.35 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 2.00 3.50 3.95 ;
        RECT  6.00 2.00 6.70 4.40 ;
        RECT  8.70 2.00 9.40 4.40 ;
        RECT  10.25 2.00 10.95 4.50 ;
        RECT  12.95 2.00 13.65 4.50 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.35 1.15 4.05 ;
        RECT  0.65 3.35 1.15 6.05 ;
        RECT  1.80 5.55 2.30 9.95 ;
        RECT  1.80 9.25 2.50 9.95 ;
        RECT  2.35 4.40 3.05 5.10 ;
        RECT  4.15 3.35 4.65 4.90 ;
        RECT  2.35 4.40 4.65 4.90 ;
        RECT  4.15 3.35 4.85 4.05 ;
        RECT  4.60 7.10 5.30 8.75 ;
        RECT  2.75 8.05 5.30 8.75 ;
        RECT  6.40 5.35 7.10 6.05 ;
        RECT  0.65 5.55 7.10 6.05 ;
        RECT  7.35 3.75 8.05 4.45 ;
        RECT  7.55 3.75 8.05 5.45 ;
        RECT  8.65 4.95 9.15 10.55 ;
        RECT  8.45 7.10 9.15 10.55 ;
        RECT  7.55 4.95 11.15 5.45 ;
        RECT  10.45 4.95 11.15 5.65 ;
        RECT  14.30 7.15 14.80 10.55 ;
        RECT  14.55 3.95 14.80 10.55 ;
        RECT  14.00 9.85 14.80 10.55 ;
        RECT  14.55 3.95 15.05 7.85 ;
        RECT  14.30 7.15 15.05 7.85 ;
        RECT  15.50 3.75 16.20 4.45 ;
        RECT  14.55 3.95 16.20 4.45 ;
    END
END NA4I1X4
MACRO NA4I2X1
    CLASS CORE ;
    FOREIGN NA4I2X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.20 3.75 10.90 4.45 ;
        RECT  10.40 3.75 10.90 8.90 ;
        RECT  10.05 7.15 10.95 8.90 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.65 6.30 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.35 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.15 7.10 3.85 11.00 ;
        RECT  4.70 9.80 5.40 11.00 ;
        RECT  6.20 7.10 6.90 11.00 ;
        RECT  11.40 7.15 12.15 11.00 ;
        RECT  14.25 7.15 14.95 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.80 ;
        RECT  3.15 2.00 3.85 3.80 ;
        RECT  6.00 2.00 6.70 4.40 ;
        RECT  8.70 2.00 9.40 4.40 ;
        RECT  11.55 2.00 12.25 4.40 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.80 7.10 1.50 10.55 ;
        RECT  1.80 3.20 2.50 3.90 ;
        RECT  2.00 3.20 2.50 7.60 ;
        RECT  0.80 7.10 2.50 7.60 ;
        RECT  2.00 4.25 4.20 4.75 ;
        RECT  3.50 4.25 4.20 4.95 ;
        RECT  4.65 3.75 5.35 4.45 ;
        RECT  4.85 3.75 5.35 8.90 ;
        RECT  4.65 7.10 5.35 8.90 ;
        RECT  6.40 5.35 7.10 6.05 ;
        RECT  4.85 5.55 7.10 6.05 ;
        RECT  7.35 3.75 8.05 4.45 ;
        RECT  7.55 3.75 8.05 5.45 ;
        RECT  7.55 4.95 9.95 5.45 ;
        RECT  8.75 4.95 9.25 10.55 ;
        RECT  8.55 7.10 9.25 10.55 ;
        RECT  8.75 4.95 9.95 5.65 ;
        RECT  12.90 7.15 13.60 7.85 ;
        RECT  13.10 3.95 13.60 10.15 ;
        RECT  12.90 9.45 13.60 10.15 ;
        RECT  13.90 3.75 14.60 4.45 ;
        RECT  13.10 3.95 14.60 4.45 ;
    END
END NA4I2X1
MACRO NA4I2X2
    CLASS CORE ;
    FOREIGN NA4I2X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.20 2.70 10.90 4.50 ;
        RECT  10.40 2.70 10.90 10.55 ;
        RECT  10.05 7.10 10.95 10.55 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.70 6.30 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.35 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.15 7.10 3.85 11.00 ;
        RECT  4.70 9.80 5.40 11.00 ;
        RECT  6.20 7.10 6.90 11.00 ;
        RECT  11.40 7.10 12.15 11.00 ;
        RECT  14.25 7.15 14.95 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.80 ;
        RECT  3.15 2.00 3.85 3.80 ;
        RECT  6.00 2.00 6.70 4.40 ;
        RECT  8.70 2.00 9.40 4.40 ;
        RECT  11.55 2.00 12.25 4.50 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.80 7.10 1.50 10.55 ;
        RECT  1.80 3.20 2.50 3.90 ;
        RECT  2.00 3.20 2.50 7.60 ;
        RECT  0.80 7.10 2.50 7.60 ;
        RECT  2.00 4.25 4.20 4.75 ;
        RECT  3.50 4.25 4.20 4.95 ;
        RECT  4.65 3.75 5.35 4.45 ;
        RECT  4.85 3.75 5.35 8.90 ;
        RECT  4.65 7.10 5.35 8.90 ;
        RECT  6.40 5.35 7.10 6.05 ;
        RECT  4.85 5.55 7.10 6.05 ;
        RECT  7.35 3.75 8.05 4.45 ;
        RECT  7.55 3.75 8.05 5.45 ;
        RECT  7.55 4.95 9.95 5.45 ;
        RECT  8.75 4.95 9.25 10.55 ;
        RECT  8.55 7.10 9.25 10.55 ;
        RECT  8.75 4.95 9.95 5.65 ;
        RECT  12.90 7.15 13.40 10.55 ;
        RECT  13.15 3.95 13.40 10.55 ;
        RECT  12.60 9.85 13.40 10.55 ;
        RECT  13.15 3.95 13.65 7.85 ;
        RECT  12.90 7.15 13.65 7.85 ;
        RECT  14.10 3.75 14.80 4.45 ;
        RECT  13.15 3.95 14.80 4.45 ;
    END
END NA4I2X2
MACRO NA4I2X4
    CLASS CORE ;
    FOREIGN NA4I2X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.60 2.70 12.35 4.50 ;
        RECT  11.85 2.70 12.35 10.55 ;
        RECT  11.45 7.10 12.35 10.55 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 14.10 6.30 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.35 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.15 7.10 3.85 11.00 ;
        RECT  4.70 9.80 5.40 11.00 ;
        RECT  6.20 7.10 6.90 11.00 ;
        RECT  10.10 7.10 10.80 11.00 ;
        RECT  12.80 7.10 13.50 11.00 ;
        RECT  15.65 7.15 16.35 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.80 ;
        RECT  3.15 2.00 3.85 3.80 ;
        RECT  6.00 2.00 6.70 4.40 ;
        RECT  8.70 2.00 9.40 4.40 ;
        RECT  10.25 2.00 10.95 4.50 ;
        RECT  12.95 2.00 13.65 4.50 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.80 7.10 1.50 10.55 ;
        RECT  1.80 3.20 2.50 3.90 ;
        RECT  2.00 3.20 2.50 7.60 ;
        RECT  0.80 7.10 2.50 7.60 ;
        RECT  2.00 4.25 4.20 4.75 ;
        RECT  3.50 4.25 4.20 4.95 ;
        RECT  4.65 3.75 5.35 4.45 ;
        RECT  4.85 3.75 5.35 8.90 ;
        RECT  4.65 7.10 5.35 8.90 ;
        RECT  6.40 5.35 7.10 6.05 ;
        RECT  4.85 5.55 7.10 6.05 ;
        RECT  7.35 3.75 8.05 4.45 ;
        RECT  7.55 3.75 8.05 5.45 ;
        RECT  8.75 4.95 9.25 10.55 ;
        RECT  8.55 7.10 9.25 10.55 ;
        RECT  7.55 4.95 11.25 5.45 ;
        RECT  10.55 4.95 11.25 5.65 ;
        RECT  14.30 7.15 14.80 10.55 ;
        RECT  14.55 3.95 14.80 10.55 ;
        RECT  14.00 9.85 14.80 10.55 ;
        RECT  14.55 3.95 15.05 7.85 ;
        RECT  14.30 7.15 15.05 7.85 ;
        RECT  15.50 3.75 16.20 4.45 ;
        RECT  14.55 3.95 16.20 4.45 ;
    END
END NA4I2X4
MACRO NA4I3X1
    CLASS CORE ;
    FOREIGN NA4I3X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.20 3.75 10.90 4.45 ;
        RECT  10.40 3.75 10.90 8.90 ;
        RECT  10.05 7.15 10.95 8.90 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.45 6.35 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.35 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.15 7.10 3.85 11.00 ;
        RECT  4.70 9.80 5.40 11.00 ;
        RECT  6.20 7.10 6.90 11.00 ;
        RECT  11.40 7.15 12.10 11.00 ;
        RECT  14.35 7.15 15.05 11.00 ;
        RECT  17.05 7.15 17.75 11.00 ;
        RECT  13.75 10.10 17.75 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.80 ;
        RECT  3.15 2.00 3.85 3.80 ;
        RECT  6.00 2.00 6.70 4.40 ;
        RECT  8.70 2.00 9.40 4.40 ;
        RECT  11.55 2.00 12.25 4.40 ;
        RECT  14.65 2.00 15.35 4.40 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.80 7.10 1.50 10.55 ;
        RECT  1.80 3.20 2.50 3.90 ;
        RECT  2.00 3.20 2.50 7.60 ;
        RECT  0.80 7.10 2.50 7.60 ;
        RECT  2.00 4.25 4.20 4.75 ;
        RECT  3.50 4.25 4.20 4.95 ;
        RECT  4.65 3.75 5.35 4.45 ;
        RECT  4.85 3.75 5.35 8.90 ;
        RECT  4.65 7.10 5.35 8.90 ;
        RECT  6.40 5.35 7.10 6.05 ;
        RECT  4.85 5.55 7.10 6.05 ;
        RECT  7.35 3.75 8.05 4.45 ;
        RECT  7.55 3.75 8.05 5.45 ;
        RECT  7.55 4.95 9.95 5.45 ;
        RECT  8.75 4.95 9.25 10.55 ;
        RECT  8.55 7.10 9.25 10.55 ;
        RECT  8.75 4.95 9.95 5.65 ;
        RECT  12.90 3.75 13.45 8.90 ;
        RECT  12.75 7.15 13.45 8.90 ;
        RECT  12.90 3.75 13.60 4.45 ;
        RECT  14.70 5.35 15.40 6.05 ;
        RECT  12.90 5.55 15.40 6.05 ;
        RECT  15.70 7.15 16.40 7.85 ;
        RECT  15.90 3.95 16.40 9.60 ;
        RECT  15.70 8.90 16.40 9.60 ;
        RECT  17.05 3.75 17.75 4.45 ;
        RECT  15.90 3.95 17.75 4.45 ;
    END
END NA4I3X1
MACRO NA4I3X2
    CLASS CORE ;
    FOREIGN NA4I3X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.20 2.70 10.90 4.50 ;
        RECT  10.40 2.70 10.90 10.55 ;
        RECT  10.05 7.15 10.95 10.55 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.45 6.35 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.35 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.15 7.10 3.85 11.00 ;
        RECT  4.70 9.80 5.40 11.00 ;
        RECT  6.20 7.10 6.90 11.00 ;
        RECT  11.40 7.10 12.10 11.00 ;
        RECT  14.35 7.15 15.05 11.00 ;
        RECT  17.05 7.15 17.75 11.00 ;
        RECT  13.85 10.10 17.75 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.80 ;
        RECT  3.15 2.00 3.85 3.80 ;
        RECT  6.00 2.00 6.70 4.40 ;
        RECT  8.70 2.00 9.40 4.40 ;
        RECT  11.55 2.00 12.25 4.50 ;
        RECT  14.70 2.00 15.40 4.40 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.80 7.10 1.50 10.55 ;
        RECT  1.80 3.20 2.50 3.90 ;
        RECT  2.00 3.20 2.50 7.60 ;
        RECT  0.80 7.10 2.50 7.60 ;
        RECT  2.00 4.25 4.20 4.75 ;
        RECT  3.50 4.25 4.20 4.95 ;
        RECT  4.65 3.75 5.35 4.45 ;
        RECT  4.85 3.75 5.35 8.90 ;
        RECT  4.65 7.10 5.35 8.90 ;
        RECT  6.40 5.35 7.10 6.05 ;
        RECT  4.85 5.55 7.10 6.05 ;
        RECT  7.35 3.75 8.05 4.45 ;
        RECT  7.55 3.75 8.05 5.45 ;
        RECT  7.55 4.95 9.95 5.45 ;
        RECT  8.75 4.95 9.25 10.55 ;
        RECT  8.55 7.10 9.25 10.55 ;
        RECT  8.75 4.95 9.95 5.65 ;
        RECT  13.05 3.75 13.55 8.90 ;
        RECT  12.85 7.10 13.55 8.90 ;
        RECT  13.05 3.75 13.75 4.45 ;
        RECT  14.70 5.35 15.40 6.05 ;
        RECT  13.05 5.55 15.40 6.05 ;
        RECT  15.70 7.15 16.40 7.85 ;
        RECT  15.90 3.95 16.40 9.60 ;
        RECT  15.70 8.90 16.40 9.60 ;
        RECT  17.05 3.75 17.75 4.45 ;
        RECT  15.90 3.95 17.75 4.45 ;
    END
END NA4I3X2
MACRO NA4I3X4
    CLASS CORE ;
    FOREIGN NA4I3X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.60 2.70 12.10 10.55 ;
        RECT  11.40 7.15 12.10 10.55 ;
        RECT  11.60 2.70 12.30 4.50 ;
        RECT  11.40 2.70 12.35 3.70 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.40 19.35 6.30 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.85 6.35 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.35 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.15 7.10 3.85 11.00 ;
        RECT  4.70 9.80 5.40 11.00 ;
        RECT  6.20 7.10 6.90 11.00 ;
        RECT  10.05 7.10 10.75 11.00 ;
        RECT  12.75 7.10 13.45 11.00 ;
        RECT  15.75 7.15 16.45 11.00 ;
        RECT  18.45 7.15 19.15 11.00 ;
        RECT  15.30 10.10 19.15 11.00 ;
        RECT  0.00 11.00 19.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.80 ;
        RECT  3.15 2.00 3.85 3.80 ;
        RECT  6.00 2.00 6.70 4.40 ;
        RECT  8.70 2.00 9.40 4.40 ;
        RECT  10.25 2.00 10.95 4.50 ;
        RECT  12.95 2.00 13.65 4.50 ;
        RECT  16.10 2.00 16.80 4.40 ;
        RECT  0.00 0.00 19.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.80 7.10 1.50 10.55 ;
        RECT  1.80 3.20 2.50 3.90 ;
        RECT  2.00 3.20 2.50 7.60 ;
        RECT  0.80 7.10 2.50 7.60 ;
        RECT  2.00 4.25 4.20 4.75 ;
        RECT  3.50 4.25 4.20 4.95 ;
        RECT  4.65 3.75 5.35 4.45 ;
        RECT  4.85 3.75 5.35 8.90 ;
        RECT  4.65 7.10 5.35 8.90 ;
        RECT  6.40 5.35 7.10 6.05 ;
        RECT  4.85 5.55 7.10 6.05 ;
        RECT  7.35 3.75 8.05 4.45 ;
        RECT  7.55 3.75 8.05 5.45 ;
        RECT  8.75 4.95 9.25 10.55 ;
        RECT  8.55 7.10 9.25 10.55 ;
        RECT  7.55 4.95 11.15 5.45 ;
        RECT  10.45 4.95 11.15 5.65 ;
        RECT  14.45 3.75 14.95 8.90 ;
        RECT  14.25 7.10 14.95 8.90 ;
        RECT  14.45 3.75 15.15 4.45 ;
        RECT  16.10 5.35 16.80 6.05 ;
        RECT  14.45 5.55 16.80 6.05 ;
        RECT  17.10 7.15 17.80 7.85 ;
        RECT  17.30 3.95 17.80 9.60 ;
        RECT  17.10 8.90 17.80 9.60 ;
        RECT  18.45 3.75 19.15 4.45 ;
        RECT  17.30 3.95 19.15 4.45 ;
    END
END NA4I3X4
MACRO NA4X1
    CLASS CORE ;
    FOREIGN NA4X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  7.40 3.75 7.90 8.90 ;
        RECT  7.40 3.75 8.10 4.45 ;
        RECT  7.25 7.15 8.15 8.90 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.40 9.85 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  0.25 6.70 1.15 7.60 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  1.65 4.10 3.05 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 9.15 1.15 11.00 ;
        RECT  0.45 10.85 2.15 11.00 ;
        RECT  3.30 7.20 4.00 11.00 ;
        RECT  8.60 7.15 9.35 11.00 ;
        RECT  7.75 10.10 9.35 11.00 ;
        RECT  11.45 7.15 12.15 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 2.00 3.50 3.65 ;
        RECT  5.50 2.00 6.20 3.65 ;
        RECT  8.75 2.00 9.45 4.40 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.05 1.15 3.75 ;
        RECT  0.65 3.05 1.15 6.05 ;
        RECT  1.80 5.55 2.30 9.85 ;
        RECT  1.80 9.15 2.50 9.85 ;
        RECT  0.65 5.55 4.45 6.05 ;
        RECT  4.15 3.00 4.85 3.70 ;
        RECT  3.75 5.55 4.45 6.25 ;
        RECT  4.35 3.00 4.85 5.00 ;
        RECT  4.35 4.50 6.95 5.00 ;
        RECT  5.85 4.50 6.35 10.55 ;
        RECT  5.65 7.15 6.35 10.55 ;
        RECT  5.85 4.50 6.95 5.20 ;
        RECT  10.10 7.15 10.80 7.85 ;
        RECT  10.30 3.95 10.80 10.55 ;
        RECT  10.10 9.85 10.80 10.55 ;
        RECT  11.10 3.75 11.80 4.45 ;
        RECT  10.30 3.95 11.80 4.45 ;
    END
END NA4X1
MACRO NA4X2
    CLASS CORE ;
    FOREIGN NA4X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  7.25 2.60 7.75 10.55 ;
        RECT  7.25 2.60 7.95 4.35 ;
        RECT  7.25 7.15 7.95 10.55 ;
        RECT  7.25 8.00 8.15 8.90 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.40 9.85 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  0.25 6.70 1.15 7.60 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  1.65 4.10 3.05 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 8.20 1.15 11.00 ;
        RECT  0.45 10.10 2.15 11.00 ;
        RECT  3.30 7.20 4.00 11.00 ;
        RECT  8.60 7.15 9.30 11.00 ;
        RECT  11.45 7.15 12.15 11.00 ;
        RECT  10.50 10.10 12.15 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 2.00 3.50 3.65 ;
        RECT  5.50 2.00 6.20 3.65 ;
        RECT  8.60 2.00 9.30 4.35 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.05 1.15 3.75 ;
        RECT  0.65 3.05 1.15 6.05 ;
        RECT  1.80 5.55 2.30 8.90 ;
        RECT  1.80 8.20 2.50 8.90 ;
        RECT  0.65 5.55 4.45 6.05 ;
        RECT  4.15 3.00 4.85 3.70 ;
        RECT  3.75 5.55 4.45 6.25 ;
        RECT  4.35 3.00 4.85 5.00 ;
        RECT  4.35 4.50 6.80 5.00 ;
        RECT  5.85 4.50 6.35 10.55 ;
        RECT  5.65 7.15 6.35 10.55 ;
        RECT  5.85 4.50 6.80 5.20 ;
        RECT  10.30 3.80 10.80 7.85 ;
        RECT  10.10 7.15 10.80 7.85 ;
        RECT  11.10 3.60 12.30 4.30 ;
        RECT  11.60 2.45 12.30 4.30 ;
        RECT  10.30 3.80 12.30 4.30 ;
    END
END NA4X2
MACRO NA4X3
    CLASS CORE ;
    FOREIGN NA4X3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  7.25 2.45 7.75 10.55 ;
        RECT  7.25 2.45 7.95 4.35 ;
        RECT  7.25 7.15 7.95 10.55 ;
        RECT  7.25 8.00 8.15 8.90 ;
        RECT  7.25 9.85 8.90 10.55 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.40 9.85 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  0.25 6.70 1.15 7.60 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  1.65 4.10 3.05 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 8.20 1.15 11.00 ;
        RECT  0.45 10.10 2.15 11.00 ;
        RECT  3.30 7.20 4.00 11.00 ;
        RECT  8.60 7.15 9.30 9.20 ;
        RECT  8.60 8.50 10.25 9.20 ;
        RECT  9.55 8.50 10.25 11.00 ;
        RECT  11.45 7.15 12.15 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 2.00 3.50 3.65 ;
        RECT  5.50 2.00 6.20 3.65 ;
        RECT  8.60 2.00 9.30 4.35 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.05 1.15 3.75 ;
        RECT  0.65 3.05 1.15 6.05 ;
        RECT  1.80 5.55 2.30 8.90 ;
        RECT  1.80 8.20 2.50 8.90 ;
        RECT  0.65 5.55 4.45 6.05 ;
        RECT  4.15 3.00 4.85 3.70 ;
        RECT  3.75 5.55 4.45 6.25 ;
        RECT  4.35 3.00 4.85 5.00 ;
        RECT  4.35 4.50 6.80 5.00 ;
        RECT  5.85 4.50 6.35 10.55 ;
        RECT  5.65 7.15 6.35 10.55 ;
        RECT  5.85 4.50 6.80 5.20 ;
        RECT  10.30 3.80 10.80 7.85 ;
        RECT  10.10 7.15 10.80 7.85 ;
        RECT  11.10 3.60 12.30 4.30 ;
        RECT  11.60 2.45 12.30 4.30 ;
        RECT  10.30 3.80 12.30 4.30 ;
    END
END NA4X3
MACRO NA4X4
    CLASS CORE ;
    FOREIGN NA4X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  7.40 2.55 7.90 10.55 ;
        RECT  7.25 7.15 7.95 10.55 ;
        RECT  7.40 2.55 8.10 4.15 ;
        RECT  7.25 8.00 8.15 8.90 ;
        RECT  7.25 9.85 9.80 10.55 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.40 9.85 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  0.25 6.70 1.15 7.60 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  1.65 9.30 2.85 10.20 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 8.20 1.15 11.00 ;
        RECT  3.30 7.20 4.00 11.00 ;
        RECT  8.60 7.20 9.30 9.20 ;
        RECT  10.45 8.60 11.15 11.00 ;
        RECT  11.45 7.20 12.15 9.20 ;
        RECT  8.60 8.60 12.15 9.20 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 2.00 3.50 4.40 ;
        RECT  5.50 2.00 6.20 4.40 ;
        RECT  8.75 2.00 9.45 4.50 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.80 1.15 4.50 ;
        RECT  0.65 3.80 1.15 5.65 ;
        RECT  0.65 5.15 2.30 5.65 ;
        RECT  1.80 5.15 2.30 8.85 ;
        RECT  1.80 8.15 2.50 8.85 ;
        RECT  4.15 3.75 4.85 4.45 ;
        RECT  3.70 5.80 4.40 6.50 ;
        RECT  1.80 6.00 4.40 6.50 ;
        RECT  4.35 3.75 4.85 5.35 ;
        RECT  4.35 4.85 6.80 5.35 ;
        RECT  5.85 4.85 6.35 10.55 ;
        RECT  5.65 7.15 6.35 10.55 ;
        RECT  5.85 4.85 6.80 5.55 ;
        RECT  10.30 3.95 10.80 7.90 ;
        RECT  10.10 7.20 10.80 7.90 ;
        RECT  11.25 3.75 11.95 4.45 ;
        RECT  11.45 2.45 11.95 4.45 ;
        RECT  10.30 3.95 11.95 4.45 ;
        RECT  11.45 2.45 12.30 3.15 ;
    END
END NA4X4
MACRO NA5I1X1
    CLASS CORE ;
    FOREIGN NA5I1X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.05 3.60 10.95 4.30 ;
        RECT  10.45 3.60 10.95 9.20 ;
        RECT  10.05 7.45 10.95 9.20 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.65 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 4.15 6.30 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.40 5.40 2.55 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.15 2.50 11.00 ;
        RECT  4.65 9.15 5.35 11.00 ;
        RECT  6.15 7.20 6.85 11.00 ;
        RECT  11.40 7.45 12.15 11.00 ;
        RECT  10.15 10.10 12.15 11.00 ;
        RECT  14.25 8.15 14.95 11.00 ;
        RECT  13.80 10.10 16.35 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.40 ;
        RECT  5.80 2.00 6.50 4.35 ;
        RECT  8.50 2.00 9.20 4.35 ;
        RECT  11.70 2.00 12.40 4.25 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.70 0.95 9.85 ;
        RECT  0.45 3.70 1.15 4.40 ;
        RECT  0.45 8.15 1.15 9.85 ;
        RECT  0.45 7.00 3.10 7.50 ;
        RECT  2.40 7.00 3.10 7.70 ;
        RECT  3.30 8.20 4.00 9.85 ;
        RECT  4.15 3.70 5.10 4.40 ;
        RECT  4.60 3.70 5.10 8.70 ;
        RECT  3.30 8.20 5.10 8.70 ;
        RECT  4.60 5.75 7.40 6.25 ;
        RECT  7.15 3.70 7.85 4.40 ;
        RECT  6.70 5.75 7.40 6.45 ;
        RECT  7.35 3.70 7.85 5.30 ;
        RECT  7.35 4.80 10.00 5.30 ;
        RECT  8.70 4.80 9.20 10.55 ;
        RECT  8.50 7.15 9.20 10.55 ;
        RECT  8.70 4.80 10.00 5.50 ;
        RECT  12.85 8.10 13.35 10.55 ;
        RECT  13.10 3.80 13.35 10.55 ;
        RECT  12.65 9.85 13.35 10.55 ;
        RECT  13.10 3.80 13.60 8.80 ;
        RECT  12.85 8.10 13.60 8.80 ;
        RECT  13.10 7.15 16.30 7.65 ;
        RECT  15.25 3.60 15.95 4.30 ;
        RECT  13.10 3.80 15.95 4.30 ;
        RECT  15.60 7.15 16.30 8.80 ;
    END
END NA5I1X1
MACRO NA5I1X2
    CLASS CORE ;
    FOREIGN NA5I1X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.45 2.55 10.95 10.55 ;
        RECT  10.05 7.10 10.95 10.55 ;
        RECT  10.40 2.55 11.10 4.30 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.65 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 4.15 6.30 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.40 5.40 2.55 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.15 2.50 11.00 ;
        RECT  4.65 9.15 5.35 11.00 ;
        RECT  6.15 7.20 6.85 11.00 ;
        RECT  11.40 7.10 12.10 11.00 ;
        RECT  14.25 8.15 14.95 11.00 ;
        RECT  13.80 10.10 16.35 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.40 ;
        RECT  5.80 2.00 6.50 4.35 ;
        RECT  8.50 2.00 9.20 4.35 ;
        RECT  11.75 2.00 12.45 4.25 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.70 0.95 9.85 ;
        RECT  0.45 3.70 1.15 4.40 ;
        RECT  0.45 8.15 1.15 9.85 ;
        RECT  0.45 7.00 3.10 7.50 ;
        RECT  2.40 7.00 3.10 7.70 ;
        RECT  3.30 8.20 4.00 9.85 ;
        RECT  4.15 3.70 5.10 4.40 ;
        RECT  4.60 3.70 5.10 8.70 ;
        RECT  3.30 8.20 5.10 8.70 ;
        RECT  4.60 5.75 7.40 6.25 ;
        RECT  7.15 3.70 7.85 4.40 ;
        RECT  6.70 5.75 7.40 6.45 ;
        RECT  7.35 3.70 7.85 5.30 ;
        RECT  7.35 4.80 10.00 5.30 ;
        RECT  8.70 4.80 9.20 10.55 ;
        RECT  8.50 7.15 9.20 10.55 ;
        RECT  8.70 4.80 10.00 5.50 ;
        RECT  12.85 8.10 13.35 10.55 ;
        RECT  13.10 3.80 13.35 10.55 ;
        RECT  12.65 9.85 13.35 10.55 ;
        RECT  13.10 3.80 13.60 8.80 ;
        RECT  12.85 8.10 13.60 8.80 ;
        RECT  13.10 7.15 16.30 7.65 ;
        RECT  15.25 3.60 15.95 4.30 ;
        RECT  13.10 3.80 15.95 4.30 ;
        RECT  15.60 7.15 16.30 8.80 ;
    END
END NA5I1X2
MACRO NA5I1X4
    CLASS CORE ;
    FOREIGN NA5I1X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.80 2.55 12.15 10.55 ;
        RECT  11.45 7.10 12.15 10.55 ;
        RECT  11.80 2.55 12.30 8.90 ;
        RECT  11.45 7.10 12.30 8.90 ;
        RECT  11.45 8.00 12.35 8.90 ;
        RECT  11.80 2.55 12.50 4.30 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 14.05 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 4.20 6.30 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.40 5.40 2.55 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.15 2.50 11.00 ;
        RECT  4.65 9.15 5.35 11.00 ;
        RECT  6.15 7.20 6.85 11.00 ;
        RECT  10.10 7.20 10.80 11.00 ;
        RECT  12.80 7.20 13.50 11.00 ;
        RECT  15.65 8.15 16.35 11.00 ;
        RECT  15.20 10.10 17.75 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.40 ;
        RECT  5.80 2.00 6.50 4.35 ;
        RECT  8.50 2.00 9.20 4.35 ;
        RECT  10.45 2.00 11.15 4.25 ;
        RECT  13.15 2.00 13.85 4.25 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.70 0.95 9.85 ;
        RECT  0.45 3.70 1.15 4.40 ;
        RECT  0.45 8.15 1.15 9.85 ;
        RECT  0.45 7.00 3.10 7.50 ;
        RECT  2.40 7.00 3.10 7.70 ;
        RECT  3.30 8.20 4.00 9.85 ;
        RECT  4.15 3.70 5.15 4.40 ;
        RECT  4.65 3.70 5.15 8.70 ;
        RECT  3.30 8.20 5.15 8.70 ;
        RECT  4.65 5.75 7.40 6.25 ;
        RECT  7.15 3.70 7.85 4.40 ;
        RECT  6.70 5.75 7.40 6.45 ;
        RECT  7.35 3.70 7.85 5.30 ;
        RECT  8.70 4.80 9.20 10.55 ;
        RECT  8.50 7.15 9.20 10.55 ;
        RECT  7.35 4.80 11.25 5.30 ;
        RECT  10.55 4.80 11.25 5.50 ;
        RECT  14.25 8.10 14.75 10.55 ;
        RECT  14.50 3.80 14.75 10.55 ;
        RECT  14.05 9.85 14.75 10.55 ;
        RECT  14.50 3.80 15.00 8.80 ;
        RECT  14.25 8.10 15.00 8.80 ;
        RECT  14.50 7.15 17.70 7.65 ;
        RECT  16.65 3.60 17.35 4.30 ;
        RECT  14.50 3.80 17.35 4.30 ;
        RECT  17.00 7.15 17.70 8.80 ;
    END
END NA5I1X4
MACRO NA5I2X1
    CLASS CORE ;
    FOREIGN NA5I2X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.45 3.75 10.95 9.20 ;
        RECT  10.05 7.45 10.95 9.20 ;
        RECT  10.45 3.75 11.25 4.45 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.35 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.65 6.45 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.35 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.15 7.10 3.85 11.00 ;
        RECT  4.70 9.80 5.40 11.00 ;
        RECT  6.20 7.10 6.90 11.00 ;
        RECT  11.40 7.45 12.15 11.00 ;
        RECT  10.20 10.10 12.15 11.00 ;
        RECT  14.25 8.15 14.95 11.00 ;
        RECT  13.80 10.10 16.35 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.80 ;
        RECT  3.15 2.00 3.85 3.80 ;
        RECT  6.00 2.00 6.70 4.40 ;
        RECT  8.70 2.00 9.40 4.40 ;
        RECT  11.90 2.00 12.60 4.40 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.80 7.10 1.50 10.55 ;
        RECT  1.80 3.20 2.50 3.90 ;
        RECT  2.00 3.20 2.50 7.60 ;
        RECT  0.80 7.10 2.50 7.60 ;
        RECT  2.00 4.25 4.20 4.75 ;
        RECT  3.50 4.25 4.20 4.95 ;
        RECT  4.65 3.75 5.35 4.45 ;
        RECT  4.85 3.75 5.35 8.90 ;
        RECT  4.65 7.10 5.35 8.90 ;
        RECT  6.40 5.35 7.10 6.05 ;
        RECT  4.85 5.55 7.10 6.05 ;
        RECT  7.35 3.75 8.05 4.45 ;
        RECT  7.55 3.75 8.05 5.45 ;
        RECT  7.55 4.95 10.00 5.45 ;
        RECT  8.75 4.95 9.25 10.55 ;
        RECT  8.55 7.10 9.25 10.55 ;
        RECT  8.75 4.95 10.00 5.65 ;
        RECT  12.85 8.10 13.35 10.55 ;
        RECT  13.10 3.95 13.35 10.55 ;
        RECT  12.65 9.85 13.35 10.55 ;
        RECT  13.10 3.95 13.60 8.80 ;
        RECT  12.85 8.10 13.60 8.80 ;
        RECT  13.10 7.15 16.30 7.65 ;
        RECT  15.25 3.75 15.95 4.45 ;
        RECT  13.10 3.95 15.95 4.45 ;
        RECT  15.60 7.15 16.30 8.80 ;
    END
END NA5I2X1
MACRO NA5I2X2
    CLASS CORE ;
    FOREIGN NA5I2X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.45 2.70 10.95 10.55 ;
        RECT  10.05 7.10 10.95 10.55 ;
        RECT  10.35 2.70 11.10 4.50 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.35 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.65 6.30 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.35 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.15 7.10 3.85 11.00 ;
        RECT  4.70 9.80 5.40 11.00 ;
        RECT  6.20 7.10 6.90 11.00 ;
        RECT  11.40 7.10 12.10 11.00 ;
        RECT  14.25 8.15 14.95 11.00 ;
        RECT  13.75 10.10 16.35 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.80 ;
        RECT  3.15 2.00 3.85 3.80 ;
        RECT  6.00 2.00 6.70 4.40 ;
        RECT  8.70 2.00 9.40 4.40 ;
        RECT  11.75 2.00 12.45 4.50 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.80 7.10 1.50 10.55 ;
        RECT  1.80 3.20 2.50 3.90 ;
        RECT  2.00 3.20 2.50 7.60 ;
        RECT  0.80 7.10 2.50 7.60 ;
        RECT  2.00 4.25 4.20 4.75 ;
        RECT  3.50 4.25 4.20 4.95 ;
        RECT  4.65 3.75 5.35 4.45 ;
        RECT  4.85 3.75 5.35 8.90 ;
        RECT  4.65 7.10 5.35 8.90 ;
        RECT  6.40 5.35 7.10 6.05 ;
        RECT  4.85 5.55 7.10 6.05 ;
        RECT  7.35 3.75 8.05 4.45 ;
        RECT  7.55 3.75 8.05 5.45 ;
        RECT  7.55 4.95 10.00 5.45 ;
        RECT  8.75 4.95 9.25 10.55 ;
        RECT  8.55 7.10 9.25 10.55 ;
        RECT  8.75 4.95 10.00 5.65 ;
        RECT  12.80 8.10 13.30 10.55 ;
        RECT  13.10 3.95 13.30 10.55 ;
        RECT  12.60 9.85 13.30 10.55 ;
        RECT  13.10 3.95 13.60 8.80 ;
        RECT  12.80 8.10 13.60 8.80 ;
        RECT  13.10 7.15 16.30 7.65 ;
        RECT  15.25 3.75 15.95 4.45 ;
        RECT  13.10 3.95 15.95 4.45 ;
        RECT  15.60 7.15 16.30 8.80 ;
    END
END NA5I2X2
MACRO NA5I2X4
    CLASS CORE ;
    FOREIGN NA5I2X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.75 2.70 12.15 10.55 ;
        RECT  11.45 7.10 12.15 10.55 ;
        RECT  11.75 2.70 12.25 8.90 ;
        RECT  11.45 7.10 12.25 8.90 ;
        RECT  11.45 8.00 12.35 8.90 ;
        RECT  11.75 2.70 12.50 4.50 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.35 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 14.05 6.30 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.35 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.15 7.10 3.85 11.00 ;
        RECT  4.70 9.80 5.40 11.00 ;
        RECT  6.20 7.10 6.90 11.00 ;
        RECT  10.10 7.10 10.80 11.00 ;
        RECT  12.80 7.10 13.50 11.00 ;
        RECT  15.65 8.15 16.35 11.00 ;
        RECT  15.15 10.10 17.75 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.80 ;
        RECT  3.15 2.00 3.85 3.80 ;
        RECT  6.00 2.00 6.70 4.40 ;
        RECT  8.70 2.00 9.40 4.40 ;
        RECT  10.40 2.00 11.10 4.50 ;
        RECT  13.15 2.00 13.85 4.50 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.80 7.10 1.50 10.55 ;
        RECT  1.80 3.20 2.50 3.90 ;
        RECT  2.00 3.20 2.50 7.60 ;
        RECT  0.80 7.10 2.50 7.60 ;
        RECT  2.00 4.25 4.20 4.75 ;
        RECT  3.50 4.25 4.20 4.95 ;
        RECT  4.65 3.75 5.35 4.45 ;
        RECT  4.85 3.75 5.35 8.90 ;
        RECT  4.65 7.10 5.35 8.90 ;
        RECT  6.40 5.35 7.10 6.05 ;
        RECT  4.85 5.55 7.10 6.05 ;
        RECT  7.35 3.75 8.05 4.45 ;
        RECT  7.55 3.75 8.05 5.45 ;
        RECT  8.75 4.95 9.25 10.55 ;
        RECT  8.55 7.10 9.25 10.55 ;
        RECT  7.55 4.95 11.25 5.45 ;
        RECT  10.55 4.95 11.25 5.65 ;
        RECT  14.20 8.10 14.70 10.55 ;
        RECT  14.50 3.95 14.70 10.55 ;
        RECT  14.00 9.85 14.70 10.55 ;
        RECT  14.50 3.95 15.00 8.80 ;
        RECT  14.20 8.10 15.00 8.80 ;
        RECT  14.50 7.15 17.70 7.65 ;
        RECT  16.65 3.75 17.35 4.45 ;
        RECT  14.50 3.95 17.35 4.45 ;
        RECT  17.00 7.15 17.70 8.80 ;
    END
END NA5I2X4
MACRO NA5I3X1
    CLASS CORE ;
    FOREIGN NA5I3X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.85 3.60 12.35 8.90 ;
        RECT  11.45 7.10 12.35 8.90 ;
        RECT  11.85 3.60 12.65 4.30 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 14.05 6.30 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.25 2.60 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.10 1.15 11.00 ;
        RECT  7.60 7.20 8.30 11.00 ;
        RECT  12.80 7.10 13.50 11.00 ;
        RECT  11.60 10.10 13.75 11.00 ;
        RECT  15.65 7.20 16.35 11.00 ;
        RECT  14.75 10.10 16.35 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.85 ;
        RECT  3.15 2.00 3.85 3.85 ;
        RECT  7.45 2.00 8.15 4.25 ;
        RECT  10.15 2.00 10.85 4.25 ;
        RECT  13.30 2.00 14.00 4.25 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.80 8.10 5.40 8.80 ;
        RECT  1.80 3.20 2.50 4.80 ;
        RECT  4.50 3.20 5.20 4.80 ;
        RECT  1.80 4.30 5.20 4.80 ;
        RECT  4.70 3.20 5.20 8.80 ;
        RECT  4.90 3.20 5.20 10.55 ;
        RECT  3.80 7.10 5.20 8.80 ;
        RECT  4.90 8.10 5.40 10.55 ;
        RECT  4.90 9.85 5.60 10.55 ;
        RECT  4.70 5.50 6.00 6.20 ;
        RECT  6.10 3.55 6.95 4.25 ;
        RECT  6.45 3.55 6.95 8.85 ;
        RECT  6.20 7.15 6.95 8.85 ;
        RECT  8.05 5.75 8.75 6.45 ;
        RECT  6.45 5.95 8.75 6.45 ;
        RECT  8.80 3.60 9.50 4.30 ;
        RECT  9.00 3.60 9.50 5.30 ;
        RECT  9.00 4.80 11.40 5.30 ;
        RECT  10.15 4.80 10.65 10.55 ;
        RECT  9.95 7.15 10.65 10.55 ;
        RECT  10.15 4.80 11.40 5.50 ;
        RECT  14.30 7.15 14.80 9.60 ;
        RECT  14.50 3.80 14.80 9.60 ;
        RECT  14.10 8.90 14.80 9.60 ;
        RECT  14.50 3.80 15.00 7.85 ;
        RECT  14.30 7.15 15.00 7.85 ;
        RECT  15.65 3.60 16.35 4.30 ;
        RECT  14.50 3.80 16.35 4.30 ;
    END
END NA5I3X1
MACRO NA5I3X2
    CLASS CORE ;
    FOREIGN NA5I3X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.85 2.55 12.35 10.55 ;
        RECT  11.45 7.10 12.35 10.55 ;
        RECT  11.80 2.55 12.50 4.30 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 14.05 6.30 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.25 2.60 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.10 1.15 11.00 ;
        RECT  7.60 7.20 8.30 11.00 ;
        RECT  12.80 7.10 13.50 11.00 ;
        RECT  15.65 7.20 16.35 11.00 ;
        RECT  14.75 10.10 16.35 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.85 ;
        RECT  3.15 2.00 3.85 3.85 ;
        RECT  7.45 2.00 8.15 4.25 ;
        RECT  10.15 2.00 10.85 4.25 ;
        RECT  13.15 2.00 13.85 4.30 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.80 8.10 5.40 8.80 ;
        RECT  1.80 3.20 2.50 4.80 ;
        RECT  4.50 3.20 5.20 4.80 ;
        RECT  1.80 4.30 5.20 4.80 ;
        RECT  4.70 3.20 5.20 8.80 ;
        RECT  4.90 3.20 5.20 10.55 ;
        RECT  3.80 7.10 5.20 8.80 ;
        RECT  4.90 8.10 5.40 10.55 ;
        RECT  4.90 9.85 5.60 10.55 ;
        RECT  4.70 5.50 6.00 6.20 ;
        RECT  6.10 3.55 6.95 4.25 ;
        RECT  6.45 3.55 6.95 8.85 ;
        RECT  6.20 7.15 6.95 8.85 ;
        RECT  8.05 5.75 8.75 6.45 ;
        RECT  6.45 5.95 8.75 6.45 ;
        RECT  8.80 3.60 9.50 4.30 ;
        RECT  9.00 3.60 9.50 5.30 ;
        RECT  9.00 4.80 11.40 5.30 ;
        RECT  10.15 4.80 10.65 10.55 ;
        RECT  9.95 7.15 10.65 10.55 ;
        RECT  10.15 4.80 11.40 5.50 ;
        RECT  14.30 7.15 14.80 9.60 ;
        RECT  14.50 3.85 14.80 9.60 ;
        RECT  14.10 8.90 14.80 9.60 ;
        RECT  14.50 3.85 15.00 7.85 ;
        RECT  14.30 7.15 15.00 7.85 ;
        RECT  15.65 3.65 16.35 4.35 ;
        RECT  14.50 3.85 16.35 4.35 ;
    END
END NA5I3X2
MACRO NA5I3X4
    CLASS CORE ;
    FOREIGN NA5I3X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  13.20 2.55 13.55 10.55 ;
        RECT  12.85 7.10 13.55 10.55 ;
        RECT  13.20 2.55 13.70 8.90 ;
        RECT  12.85 7.10 13.70 8.90 ;
        RECT  12.85 8.00 13.75 8.90 ;
        RECT  13.20 2.55 13.90 4.30 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.45 6.30 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.25 2.60 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.10 1.15 11.00 ;
        RECT  7.60 7.20 8.30 11.00 ;
        RECT  11.50 7.10 12.20 11.00 ;
        RECT  14.20 7.10 14.90 11.00 ;
        RECT  17.05 7.20 17.75 11.00 ;
        RECT  16.15 10.10 17.75 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.85 ;
        RECT  3.15 2.00 3.85 3.85 ;
        RECT  7.45 2.00 8.15 4.25 ;
        RECT  10.15 2.00 10.85 4.25 ;
        RECT  11.85 2.00 12.55 4.30 ;
        RECT  14.55 2.00 15.25 4.30 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.80 8.10 5.40 8.80 ;
        RECT  1.80 3.20 2.50 4.80 ;
        RECT  4.50 3.20 5.20 4.80 ;
        RECT  1.80 4.30 5.20 4.80 ;
        RECT  4.70 3.20 5.20 8.80 ;
        RECT  4.90 3.20 5.20 10.55 ;
        RECT  3.80 7.10 5.20 8.80 ;
        RECT  4.90 8.10 5.40 10.55 ;
        RECT  4.90 9.85 5.60 10.55 ;
        RECT  4.70 5.50 6.00 6.20 ;
        RECT  6.10 3.55 6.95 4.25 ;
        RECT  6.45 3.55 6.95 8.85 ;
        RECT  6.20 7.15 6.95 8.85 ;
        RECT  8.05 5.75 8.75 6.45 ;
        RECT  6.45 5.95 8.75 6.45 ;
        RECT  8.80 3.60 9.50 4.30 ;
        RECT  9.00 3.60 9.50 5.30 ;
        RECT  10.15 4.80 10.65 10.55 ;
        RECT  9.95 7.15 10.65 10.55 ;
        RECT  9.00 4.80 12.65 5.30 ;
        RECT  11.95 4.80 12.65 5.50 ;
        RECT  15.70 7.15 16.20 9.60 ;
        RECT  15.90 3.85 16.20 9.60 ;
        RECT  15.50 8.90 16.20 9.60 ;
        RECT  15.90 3.85 16.40 7.85 ;
        RECT  15.70 7.15 16.40 7.85 ;
        RECT  17.05 3.65 17.75 4.35 ;
        RECT  15.90 3.85 17.75 4.35 ;
    END
END NA5I3X4
MACRO NA5I4X1
    CLASS CORE ;
    FOREIGN NA5I4X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.85 3.75 12.10 8.90 ;
        RECT  11.40 5.40 12.10 8.90 ;
        RECT  11.85 3.75 12.35 6.30 ;
        RECT  11.40 5.40 12.35 6.30 ;
        RECT  11.85 3.75 12.60 4.45 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END E
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.40 19.35 6.30 ;
        END
    END DN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.25 2.60 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.10 1.15 11.00 ;
        RECT  7.55 7.10 8.25 11.00 ;
        RECT  12.75 7.10 13.45 11.00 ;
        RECT  11.60 10.10 13.75 11.00 ;
        RECT  15.60 7.15 16.30 11.00 ;
        RECT  18.45 7.10 19.15 11.00 ;
        RECT  14.70 10.10 19.15 11.00 ;
        RECT  0.00 11.00 19.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.85 ;
        RECT  3.15 2.00 3.85 3.85 ;
        RECT  7.45 2.00 8.15 4.40 ;
        RECT  10.15 2.00 10.85 4.40 ;
        RECT  13.25 2.00 13.95 4.40 ;
        RECT  18.45 2.00 19.15 4.45 ;
        RECT  0.00 0.00 19.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.80 8.10 5.40 8.80 ;
        RECT  1.80 3.20 2.50 4.80 ;
        RECT  4.50 3.20 5.20 4.80 ;
        RECT  1.80 4.30 5.20 4.80 ;
        RECT  4.70 3.20 5.20 8.80 ;
        RECT  4.90 3.20 5.20 10.55 ;
        RECT  3.80 7.10 5.20 8.80 ;
        RECT  4.90 8.10 5.40 10.55 ;
        RECT  4.90 9.85 5.60 10.55 ;
        RECT  4.70 5.50 6.00 6.20 ;
        RECT  6.10 3.75 6.95 4.45 ;
        RECT  6.45 3.75 6.95 8.90 ;
        RECT  6.20 7.10 6.95 8.90 ;
        RECT  8.00 5.75 8.70 6.45 ;
        RECT  6.45 5.95 8.70 6.45 ;
        RECT  8.80 3.75 9.50 4.45 ;
        RECT  9.00 3.75 9.50 5.35 ;
        RECT  9.00 4.85 10.60 5.35 ;
        RECT  10.10 4.85 10.60 10.55 ;
        RECT  9.90 7.15 10.60 10.55 ;
        RECT  10.10 5.75 10.95 6.45 ;
        RECT  14.25 7.15 14.80 9.60 ;
        RECT  14.45 3.95 14.80 9.60 ;
        RECT  14.10 8.90 14.80 9.60 ;
        RECT  14.45 3.95 14.95 7.85 ;
        RECT  14.25 7.15 14.95 7.85 ;
        RECT  15.60 3.75 16.30 4.45 ;
        RECT  14.45 3.95 16.30 4.45 ;
        RECT  15.95 2.60 16.65 3.30 ;
        RECT  15.95 2.80 17.60 3.30 ;
        RECT  17.10 2.80 17.60 8.90 ;
        RECT  17.10 3.75 17.80 4.45 ;
        RECT  17.10 7.10 17.80 8.90 ;
    END
END NA5I4X1
MACRO NA5I4X2
    CLASS CORE ;
    FOREIGN NA5I4X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.65 2.70 12.10 10.55 ;
        RECT  11.40 5.40 12.10 10.55 ;
        RECT  11.65 2.70 12.35 6.30 ;
        RECT  11.40 5.40 12.35 6.30 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END E
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.40 19.35 6.30 ;
        END
    END DN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.25 2.60 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.10 1.15 11.00 ;
        RECT  7.55 7.10 8.25 11.00 ;
        RECT  12.75 7.10 13.45 11.00 ;
        RECT  15.60 7.15 16.30 11.00 ;
        RECT  18.45 7.10 19.15 11.00 ;
        RECT  14.70 10.10 19.15 11.00 ;
        RECT  0.00 11.00 19.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.85 ;
        RECT  3.15 2.00 3.85 3.85 ;
        RECT  7.45 2.00 8.15 4.40 ;
        RECT  10.15 2.00 10.85 4.40 ;
        RECT  13.00 2.00 13.70 4.50 ;
        RECT  18.45 2.00 19.15 4.45 ;
        RECT  0.00 0.00 19.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.80 8.10 5.40 8.80 ;
        RECT  1.80 3.20 2.50 4.80 ;
        RECT  4.50 3.20 5.20 4.80 ;
        RECT  1.80 4.30 5.20 4.80 ;
        RECT  4.70 3.20 5.20 8.80 ;
        RECT  4.90 3.20 5.20 10.55 ;
        RECT  3.80 7.10 5.20 8.80 ;
        RECT  4.90 8.10 5.40 10.55 ;
        RECT  4.90 9.85 5.60 10.55 ;
        RECT  4.70 5.50 6.00 6.20 ;
        RECT  6.10 3.75 6.95 4.45 ;
        RECT  6.45 3.75 6.95 8.90 ;
        RECT  6.20 7.10 6.95 8.90 ;
        RECT  8.00 5.75 8.70 6.45 ;
        RECT  6.45 5.95 8.70 6.45 ;
        RECT  8.80 3.75 9.50 4.45 ;
        RECT  9.00 3.75 9.50 5.35 ;
        RECT  9.00 4.85 10.60 5.35 ;
        RECT  10.10 4.85 10.60 10.55 ;
        RECT  9.90 7.15 10.60 10.55 ;
        RECT  10.10 5.75 10.95 6.45 ;
        RECT  14.25 7.15 14.80 9.60 ;
        RECT  14.45 3.95 14.80 9.60 ;
        RECT  14.10 8.90 14.80 9.60 ;
        RECT  14.45 3.95 14.95 7.85 ;
        RECT  14.25 7.15 14.95 7.85 ;
        RECT  15.60 3.75 16.30 4.45 ;
        RECT  14.45 3.95 16.30 4.45 ;
        RECT  15.95 2.60 16.65 3.30 ;
        RECT  15.95 2.80 17.60 3.30 ;
        RECT  17.10 2.80 17.60 8.90 ;
        RECT  17.10 3.75 17.80 4.45 ;
        RECT  17.10 7.10 17.80 8.90 ;
    END
END NA5I4X2
MACRO NA5I4X4
    CLASS CORE ;
    FOREIGN NA5I4X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  13.05 2.70 13.50 10.55 ;
        RECT  12.80 5.40 13.50 10.55 ;
        RECT  13.05 2.70 13.75 6.30 ;
        RECT  12.80 5.40 13.75 6.30 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END E
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END DN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.25 2.60 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.10 1.15 11.00 ;
        RECT  7.55 7.10 8.25 11.00 ;
        RECT  11.45 7.10 12.15 11.00 ;
        RECT  14.15 7.10 14.85 11.00 ;
        RECT  17.00 7.15 17.70 11.00 ;
        RECT  19.85 7.10 20.55 11.00 ;
        RECT  16.10 10.10 20.55 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.85 ;
        RECT  3.15 2.00 3.85 3.85 ;
        RECT  7.45 2.00 8.15 4.40 ;
        RECT  10.15 2.00 10.85 4.40 ;
        RECT  11.70 2.00 12.40 4.50 ;
        RECT  14.40 2.00 15.10 4.50 ;
        RECT  19.85 2.00 20.55 4.45 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.80 8.10 5.40 8.80 ;
        RECT  1.80 3.20 2.50 4.80 ;
        RECT  4.50 3.20 5.20 4.80 ;
        RECT  1.80 4.30 5.20 4.80 ;
        RECT  4.70 3.20 5.20 8.80 ;
        RECT  4.90 3.20 5.20 10.55 ;
        RECT  3.80 7.10 5.20 8.80 ;
        RECT  4.90 8.10 5.40 10.55 ;
        RECT  4.90 9.85 5.60 10.55 ;
        RECT  4.70 5.50 6.00 6.20 ;
        RECT  6.10 3.75 6.95 4.45 ;
        RECT  6.45 3.75 6.95 8.90 ;
        RECT  6.20 7.10 6.95 8.90 ;
        RECT  8.00 5.75 8.70 6.45 ;
        RECT  6.45 5.95 8.70 6.45 ;
        RECT  8.80 3.75 9.50 4.45 ;
        RECT  9.00 3.75 9.50 5.35 ;
        RECT  9.00 4.85 10.60 5.35 ;
        RECT  10.10 4.85 10.60 10.55 ;
        RECT  9.90 7.15 10.60 10.55 ;
        RECT  10.10 5.95 12.35 6.45 ;
        RECT  11.65 5.95 12.35 6.65 ;
        RECT  15.65 7.15 16.20 9.60 ;
        RECT  15.85 3.95 16.20 9.60 ;
        RECT  15.50 8.90 16.20 9.60 ;
        RECT  15.85 3.95 16.35 7.85 ;
        RECT  15.65 7.15 16.35 7.85 ;
        RECT  17.00 3.75 17.70 4.45 ;
        RECT  15.85 3.95 17.70 4.45 ;
        RECT  17.35 2.60 18.05 3.30 ;
        RECT  17.35 2.80 19.00 3.30 ;
        RECT  18.50 2.80 19.00 8.90 ;
        RECT  18.50 3.75 19.20 4.45 ;
        RECT  18.50 7.10 19.20 8.90 ;
    END
END NA5I4X4
MACRO NA5X1
    CLASS CORE ;
    FOREIGN NA5X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.80 3.75 9.30 8.90 ;
        RECT  8.80 3.75 9.50 4.45 ;
        RECT  8.65 7.15 9.55 8.90 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 11.25 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  0.25 6.70 1.15 7.60 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.55 7.60 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 4.45 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 9.15 2.55 11.00 ;
        RECT  4.70 7.20 5.40 11.00 ;
        RECT  10.00 7.15 10.75 11.00 ;
        RECT  9.15 10.10 10.75 11.00 ;
        RECT  12.85 7.15 13.55 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  4.20 2.00 4.90 3.65 ;
        RECT  6.90 2.00 7.60 3.65 ;
        RECT  10.15 2.00 10.85 4.40 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.85 2.80 1.55 3.50 ;
        RECT  0.50 8.20 1.20 9.85 ;
        RECT  1.05 2.80 1.55 6.05 ;
        RECT  0.50 8.20 3.90 8.70 ;
        RECT  3.40 5.55 3.90 9.85 ;
        RECT  3.20 8.20 3.90 9.85 ;
        RECT  1.05 5.55 5.85 6.05 ;
        RECT  5.55 3.00 6.25 3.70 ;
        RECT  5.15 5.55 5.85 6.25 ;
        RECT  5.75 3.00 6.25 5.00 ;
        RECT  5.75 4.50 8.35 5.00 ;
        RECT  7.25 4.50 7.75 10.55 ;
        RECT  7.05 7.15 7.75 10.55 ;
        RECT  7.25 4.50 8.35 5.20 ;
        RECT  11.50 7.15 12.20 7.85 ;
        RECT  11.70 3.95 12.20 10.55 ;
        RECT  11.50 9.85 12.20 10.55 ;
        RECT  12.50 3.75 13.20 4.45 ;
        RECT  11.70 3.95 13.20 4.45 ;
    END
END NA5X1
MACRO NA5X2
    CLASS CORE ;
    FOREIGN NA5X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.65 2.60 9.15 10.55 ;
        RECT  8.65 2.60 9.35 4.35 ;
        RECT  8.65 7.15 9.35 10.55 ;
        RECT  8.65 8.00 9.55 8.90 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 11.25 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  0.25 6.70 1.15 7.60 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.55 7.60 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 4.45 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 9.05 2.55 11.00 ;
        RECT  4.70 7.20 5.40 11.00 ;
        RECT  10.00 7.15 10.70 11.00 ;
        RECT  12.85 7.15 13.55 11.00 ;
        RECT  11.90 10.10 13.55 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  4.20 2.00 4.90 3.65 ;
        RECT  6.90 2.00 7.60 3.65 ;
        RECT  10.00 2.00 10.70 4.35 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.85 2.80 1.55 3.50 ;
        RECT  0.70 8.10 1.20 9.75 ;
        RECT  0.50 9.05 1.20 9.75 ;
        RECT  1.05 2.80 1.55 6.05 ;
        RECT  0.70 8.10 3.70 8.60 ;
        RECT  3.20 5.55 3.70 9.75 ;
        RECT  3.20 9.05 3.90 9.75 ;
        RECT  1.05 5.55 5.85 6.05 ;
        RECT  5.55 3.00 6.25 3.70 ;
        RECT  5.15 5.55 5.85 6.25 ;
        RECT  5.75 3.00 6.25 5.00 ;
        RECT  5.75 4.50 8.20 5.00 ;
        RECT  7.25 4.50 7.75 10.55 ;
        RECT  7.05 7.15 7.75 10.55 ;
        RECT  7.25 4.50 8.20 5.20 ;
        RECT  11.70 3.80 12.20 7.85 ;
        RECT  11.50 7.15 12.20 7.85 ;
        RECT  12.50 3.60 13.70 4.30 ;
        RECT  13.00 2.45 13.70 4.30 ;
        RECT  11.70 3.80 13.70 4.30 ;
    END
END NA5X2
MACRO NA5X3
    CLASS CORE ;
    FOREIGN NA5X3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.65 2.45 9.15 10.55 ;
        RECT  8.65 2.45 9.35 4.35 ;
        RECT  8.65 7.15 9.35 10.55 ;
        RECT  8.65 8.00 9.55 8.90 ;
        RECT  8.65 9.85 10.30 10.55 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 11.25 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  0.25 6.70 1.15 7.60 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.55 7.60 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 4.45 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 9.00 2.55 11.00 ;
        RECT  4.70 7.20 5.40 11.00 ;
        RECT  10.00 7.15 10.70 9.20 ;
        RECT  10.00 8.50 11.65 9.20 ;
        RECT  10.95 8.50 11.65 11.00 ;
        RECT  12.85 7.15 13.55 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  4.20 2.00 4.90 3.65 ;
        RECT  6.90 2.00 7.60 3.65 ;
        RECT  10.00 2.00 10.70 4.35 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.85 3.05 1.55 3.75 ;
        RECT  0.70 8.05 1.20 9.70 ;
        RECT  0.50 9.00 1.20 9.70 ;
        RECT  1.05 3.05 1.55 6.05 ;
        RECT  0.70 8.05 3.70 8.55 ;
        RECT  3.20 5.55 3.70 9.70 ;
        RECT  3.20 9.00 3.90 9.70 ;
        RECT  1.05 5.55 5.85 6.05 ;
        RECT  5.55 3.00 6.25 3.70 ;
        RECT  5.15 5.55 5.85 6.25 ;
        RECT  5.75 3.00 6.25 5.00 ;
        RECT  5.75 4.50 8.20 5.00 ;
        RECT  7.25 4.50 7.75 10.55 ;
        RECT  7.05 7.15 7.75 10.55 ;
        RECT  7.25 4.50 8.20 5.20 ;
        RECT  11.70 3.80 12.20 7.85 ;
        RECT  11.50 7.15 12.20 7.85 ;
        RECT  12.50 3.60 13.70 4.30 ;
        RECT  13.00 2.45 13.70 4.30 ;
        RECT  11.70 3.80 13.70 4.30 ;
    END
END NA5X3
MACRO NA5X4
    CLASS CORE ;
    FOREIGN NA5X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.80 2.55 9.30 10.55 ;
        RECT  8.65 7.15 9.35 10.55 ;
        RECT  8.80 2.55 9.50 4.15 ;
        RECT  8.65 8.00 9.55 8.90 ;
        RECT  8.65 9.85 11.20 10.55 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 11.25 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  0.25 6.70 1.15 7.60 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.55 7.60 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 4.25 7.60 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 9.00 2.55 11.00 ;
        RECT  4.70 9.00 5.40 11.00 ;
        RECT  10.00 7.20 10.70 9.20 ;
        RECT  11.85 8.60 12.55 11.00 ;
        RECT  12.85 7.20 13.55 9.20 ;
        RECT  10.00 8.60 13.55 9.20 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  4.20 2.00 4.90 4.40 ;
        RECT  6.90 2.00 7.60 4.40 ;
        RECT  10.15 2.00 10.85 4.50 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.85 3.50 1.55 4.20 ;
        RECT  0.70 8.05 1.20 9.60 ;
        RECT  0.50 8.90 1.20 9.60 ;
        RECT  1.05 3.50 1.55 5.65 ;
        RECT  3.20 8.05 3.90 9.60 ;
        RECT  1.05 5.15 5.20 5.65 ;
        RECT  4.70 5.15 5.20 8.55 ;
        RECT  0.70 8.05 5.20 8.55 ;
        RECT  5.55 3.75 6.25 4.45 ;
        RECT  4.70 5.80 5.80 6.50 ;
        RECT  5.75 3.75 6.25 5.35 ;
        RECT  5.75 4.85 8.20 5.35 ;
        RECT  7.25 4.85 7.75 10.55 ;
        RECT  7.05 8.05 7.75 10.55 ;
        RECT  7.25 4.85 8.20 5.55 ;
        RECT  11.70 3.95 12.20 7.90 ;
        RECT  11.50 7.20 12.20 7.90 ;
        RECT  12.65 3.75 13.35 4.45 ;
        RECT  12.85 2.45 13.35 4.45 ;
        RECT  11.70 3.95 13.35 4.45 ;
        RECT  12.85 2.45 13.70 3.15 ;
    END
END NA5X4
MACRO NA6I1X1
    CLASS CORE ;
    FOREIGN NA6I1X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.85 3.65 12.35 8.90 ;
        RECT  11.45 7.15 12.35 8.90 ;
        RECT  11.85 3.65 12.65 4.35 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 14.05 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.40 7.60 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 4.15 6.30 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.40 5.40 2.55 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.15 2.50 11.00 ;
        RECT  4.65 9.15 5.35 11.00 ;
        RECT  7.50 7.20 8.20 11.00 ;
        RECT  12.80 7.15 13.55 11.00 ;
        RECT  11.50 10.10 13.55 11.00 ;
        RECT  15.65 7.75 16.35 11.00 ;
        RECT  15.20 10.10 17.75 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.40 ;
        RECT  7.00 2.00 7.70 4.35 ;
        RECT  9.70 2.00 10.40 4.35 ;
        RECT  13.30 2.00 14.00 4.30 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.70 0.95 9.85 ;
        RECT  0.45 3.70 1.15 4.40 ;
        RECT  0.45 8.15 1.15 9.85 ;
        RECT  0.45 7.00 3.10 7.50 ;
        RECT  2.40 7.00 3.10 7.70 ;
        RECT  3.30 8.20 4.00 9.85 ;
        RECT  5.15 3.50 5.85 4.20 ;
        RECT  5.35 3.50 5.85 6.25 ;
        RECT  3.30 8.20 6.70 8.70 ;
        RECT  6.20 5.75 6.70 9.85 ;
        RECT  6.00 8.20 6.70 9.85 ;
        RECT  5.35 5.75 8.65 6.25 ;
        RECT  8.35 3.70 9.05 4.40 ;
        RECT  7.95 5.75 8.65 6.45 ;
        RECT  8.55 3.70 9.05 5.30 ;
        RECT  8.55 4.80 11.40 5.30 ;
        RECT  10.05 4.80 10.55 10.55 ;
        RECT  9.85 7.15 10.55 10.55 ;
        RECT  10.05 4.80 11.40 5.50 ;
        RECT  14.25 7.70 14.75 10.15 ;
        RECT  14.50 3.85 14.75 10.15 ;
        RECT  14.05 9.45 14.75 10.15 ;
        RECT  14.50 3.85 15.00 8.40 ;
        RECT  14.25 7.70 15.00 8.40 ;
        RECT  14.50 6.75 17.70 7.25 ;
        RECT  16.65 3.65 17.35 4.35 ;
        RECT  14.50 3.85 17.35 4.35 ;
        RECT  17.00 6.75 17.70 8.40 ;
    END
END NA6I1X1
MACRO NA6I1X2
    CLASS CORE ;
    FOREIGN NA6I1X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.85 2.70 12.15 10.55 ;
        RECT  11.45 7.15 12.15 10.55 ;
        RECT  11.85 2.70 12.35 8.90 ;
        RECT  11.45 7.15 12.35 8.90 ;
        RECT  11.80 2.70 12.50 4.30 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 14.05 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.40 7.60 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 4.15 6.30 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.40 5.40 2.55 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.15 2.50 11.00 ;
        RECT  4.65 9.15 5.35 11.00 ;
        RECT  7.50 7.15 8.20 11.00 ;
        RECT  12.80 7.15 13.50 11.00 ;
        RECT  15.65 7.75 16.35 11.00 ;
        RECT  15.20 10.10 17.75 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.40 ;
        RECT  7.00 2.00 7.70 4.35 ;
        RECT  9.70 2.00 10.40 4.35 ;
        RECT  13.15 2.00 13.85 4.30 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.70 0.95 9.85 ;
        RECT  0.45 3.70 1.15 4.40 ;
        RECT  0.45 8.15 1.15 9.85 ;
        RECT  0.45 7.00 3.10 7.50 ;
        RECT  2.40 7.00 3.10 7.70 ;
        RECT  3.30 8.20 4.00 9.85 ;
        RECT  5.15 3.50 5.85 4.20 ;
        RECT  5.35 3.50 5.85 6.25 ;
        RECT  3.30 8.20 6.70 8.70 ;
        RECT  6.20 5.75 6.70 9.85 ;
        RECT  6.00 8.20 6.70 9.85 ;
        RECT  5.35 5.75 8.65 6.25 ;
        RECT  8.35 3.70 9.05 4.40 ;
        RECT  7.95 5.75 8.65 6.45 ;
        RECT  8.55 3.70 9.05 5.30 ;
        RECT  8.55 4.80 11.40 5.30 ;
        RECT  10.05 4.80 10.55 10.55 ;
        RECT  9.85 7.15 10.55 10.55 ;
        RECT  10.05 4.80 11.40 5.50 ;
        RECT  14.25 7.70 14.75 10.15 ;
        RECT  14.50 3.80 14.75 10.15 ;
        RECT  14.05 9.45 14.75 10.15 ;
        RECT  14.50 3.80 15.00 8.40 ;
        RECT  14.25 7.70 15.00 8.40 ;
        RECT  14.50 6.75 17.70 7.25 ;
        RECT  16.65 3.60 17.35 4.30 ;
        RECT  14.50 3.80 17.35 4.30 ;
        RECT  17.00 6.75 17.70 8.40 ;
    END
END NA6I1X2
MACRO NA6I1X4
    CLASS CORE ;
    FOREIGN NA6I1X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  13.20 2.70 13.55 10.55 ;
        RECT  12.85 7.15 13.55 10.55 ;
        RECT  13.20 2.70 13.70 8.90 ;
        RECT  12.85 7.15 13.70 8.90 ;
        RECT  12.85 8.00 13.75 8.90 ;
        RECT  13.20 2.70 13.90 4.30 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.40 19.35 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.45 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.40 7.60 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 4.15 6.30 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.40 5.40 2.55 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.15 2.50 11.00 ;
        RECT  4.65 9.15 5.35 11.00 ;
        RECT  7.50 7.15 8.20 11.00 ;
        RECT  11.50 7.15 12.20 11.00 ;
        RECT  14.20 7.15 14.90 11.00 ;
        RECT  17.05 7.75 17.75 11.00 ;
        RECT  16.60 10.10 19.15 11.00 ;
        RECT  0.00 11.00 19.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.40 ;
        RECT  7.00 2.00 7.70 4.35 ;
        RECT  9.70 2.00 10.40 4.35 ;
        RECT  11.85 2.00 12.55 4.30 ;
        RECT  14.55 2.00 15.25 4.30 ;
        RECT  0.00 0.00 19.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 3.70 0.95 9.85 ;
        RECT  0.45 3.70 1.15 4.40 ;
        RECT  0.45 8.15 1.15 9.85 ;
        RECT  0.45 7.00 3.10 7.50 ;
        RECT  2.40 7.00 3.10 7.70 ;
        RECT  3.30 8.20 4.00 9.85 ;
        RECT  5.15 3.50 5.85 4.20 ;
        RECT  5.35 3.50 5.85 6.25 ;
        RECT  3.30 8.20 6.70 8.70 ;
        RECT  6.20 5.75 6.70 9.85 ;
        RECT  6.00 8.20 6.70 9.85 ;
        RECT  5.35 5.75 8.65 6.25 ;
        RECT  8.35 3.70 9.05 4.40 ;
        RECT  7.95 5.75 8.65 6.45 ;
        RECT  8.55 3.70 9.05 5.30 ;
        RECT  10.05 4.80 10.55 10.55 ;
        RECT  9.85 7.15 10.55 10.55 ;
        RECT  8.55 4.80 12.65 5.30 ;
        RECT  11.95 4.80 12.65 5.50 ;
        RECT  15.65 7.70 16.15 10.15 ;
        RECT  15.90 3.80 16.15 10.15 ;
        RECT  15.45 9.45 16.15 10.15 ;
        RECT  15.90 3.80 16.40 8.40 ;
        RECT  15.65 7.70 16.40 8.40 ;
        RECT  15.90 6.75 19.10 7.25 ;
        RECT  18.05 3.60 18.75 4.30 ;
        RECT  15.90 3.80 18.75 4.30 ;
        RECT  18.40 6.75 19.10 8.40 ;
    END
END NA6I1X4
MACRO NA6I2X1
    CLASS CORE ;
    FOREIGN NA6I2X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  13.25 3.60 13.75 8.90 ;
        RECT  12.85 7.15 13.75 8.90 ;
        RECT  13.25 3.60 14.05 4.30 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.40 19.35 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.45 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.40 6.30 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  8.55 5.40 9.55 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.40 5.40 2.55 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.15 2.50 11.00 ;
        RECT  4.65 9.15 5.35 11.00 ;
        RECT  9.00 7.20 9.70 11.00 ;
        RECT  14.20 7.15 14.95 11.00 ;
        RECT  13.00 10.10 14.95 11.00 ;
        RECT  17.05 7.75 17.75 11.00 ;
        RECT  16.65 10.10 19.15 11.00 ;
        RECT  0.00 11.00 19.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.40 ;
        RECT  8.85 2.00 9.55 4.35 ;
        RECT  11.55 2.00 12.25 4.35 ;
        RECT  14.70 2.00 15.40 4.25 ;
        RECT  0.00 0.00 19.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.30 7.15 8.20 7.50 ;
        RECT  0.45 3.70 0.95 9.85 ;
        RECT  0.45 3.70 1.15 4.40 ;
        RECT  0.45 8.15 1.15 9.85 ;
        RECT  0.45 7.00 2.85 7.50 ;
        RECT  2.15 7.00 2.85 7.70 ;
        RECT  3.30 3.70 3.80 9.85 ;
        RECT  3.30 8.20 4.00 9.85 ;
        RECT  4.30 7.00 5.00 7.70 ;
        RECT  5.15 2.65 5.85 4.20 ;
        RECT  3.30 3.70 5.85 4.20 ;
        RECT  3.30 8.20 6.50 8.70 ;
        RECT  6.00 8.20 6.50 9.85 ;
        RECT  6.00 9.15 6.70 9.85 ;
        RECT  7.15 2.45 7.85 3.15 ;
        RECT  5.15 2.65 7.85 3.15 ;
        RECT  7.50 3.65 8.00 8.85 ;
        RECT  4.30 7.00 8.00 7.50 ;
        RECT  7.50 3.65 8.20 4.35 ;
        RECT  7.50 7.15 8.20 8.85 ;
        RECT  10.20 3.70 10.90 4.40 ;
        RECT  10.40 3.70 10.90 5.30 ;
        RECT  10.40 4.80 12.80 5.30 ;
        RECT  11.55 4.80 12.05 10.55 ;
        RECT  11.35 7.15 12.05 10.55 ;
        RECT  11.55 4.80 12.80 5.50 ;
        RECT  15.70 7.70 16.20 10.55 ;
        RECT  15.90 3.80 16.20 10.55 ;
        RECT  15.50 9.85 16.20 10.55 ;
        RECT  15.90 3.80 16.40 8.40 ;
        RECT  15.70 7.70 16.40 8.40 ;
        RECT  15.90 6.75 19.10 7.25 ;
        RECT  18.05 3.60 18.75 4.30 ;
        RECT  15.90 3.80 18.75 4.30 ;
        RECT  18.40 6.75 19.10 8.40 ;
    END
END NA6I2X1
MACRO NA6I2X2
    CLASS CORE ;
    FOREIGN NA6I2X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  13.20 2.60 13.55 10.55 ;
        RECT  12.85 7.15 13.55 10.55 ;
        RECT  13.20 2.60 13.70 8.90 ;
        RECT  12.85 7.15 13.70 8.90 ;
        RECT  12.85 8.00 13.75 8.90 ;
        RECT  13.20 2.60 13.90 4.30 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.40 19.35 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.45 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.40 6.30 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  8.55 5.40 9.55 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.40 5.40 2.55 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.15 2.50 11.00 ;
        RECT  4.65 9.15 5.35 11.00 ;
        RECT  9.00 7.20 9.70 11.00 ;
        RECT  14.20 7.20 14.90 11.00 ;
        RECT  17.05 7.75 17.75 11.00 ;
        RECT  16.65 10.10 19.15 11.00 ;
        RECT  0.00 11.00 19.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.40 ;
        RECT  8.85 2.00 9.55 4.35 ;
        RECT  11.55 2.00 12.25 4.35 ;
        RECT  14.55 2.00 15.25 4.30 ;
        RECT  0.00 0.00 19.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.30 7.15 8.20 7.50 ;
        RECT  0.45 3.70 0.95 9.85 ;
        RECT  0.45 3.70 1.15 4.40 ;
        RECT  0.45 8.15 1.15 9.85 ;
        RECT  0.45 7.00 2.85 7.50 ;
        RECT  2.15 7.00 2.85 7.70 ;
        RECT  3.30 3.70 3.80 9.85 ;
        RECT  3.30 8.20 4.00 9.85 ;
        RECT  4.30 7.00 5.00 7.70 ;
        RECT  5.15 2.65 5.85 4.20 ;
        RECT  3.30 3.70 5.85 4.20 ;
        RECT  3.30 8.20 6.50 8.70 ;
        RECT  6.00 8.20 6.50 9.85 ;
        RECT  6.00 9.15 6.70 9.85 ;
        RECT  7.15 2.45 7.85 3.15 ;
        RECT  5.15 2.65 7.85 3.15 ;
        RECT  7.50 3.65 8.00 8.85 ;
        RECT  4.30 7.00 8.00 7.50 ;
        RECT  7.50 3.65 8.20 4.35 ;
        RECT  7.50 7.15 8.20 8.85 ;
        RECT  10.20 3.70 10.90 4.40 ;
        RECT  10.40 3.70 10.90 5.30 ;
        RECT  10.40 4.80 12.75 5.30 ;
        RECT  11.55 4.80 12.05 10.55 ;
        RECT  11.35 7.15 12.05 10.55 ;
        RECT  11.55 4.80 12.75 5.50 ;
        RECT  15.70 7.70 16.20 10.55 ;
        RECT  15.90 3.80 16.20 10.55 ;
        RECT  15.50 9.85 16.20 10.55 ;
        RECT  15.90 3.80 16.40 8.40 ;
        RECT  15.70 7.70 16.40 8.40 ;
        RECT  15.90 6.75 19.10 7.25 ;
        RECT  18.05 3.60 18.75 4.30 ;
        RECT  15.90 3.80 18.75 4.30 ;
        RECT  18.40 6.75 19.10 8.40 ;
    END
END NA6I2X2
MACRO NA6I2X4
    CLASS CORE ;
    FOREIGN NA6I2X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  14.60 2.60 14.95 10.55 ;
        RECT  14.25 7.15 14.95 10.55 ;
        RECT  14.60 2.60 15.10 8.90 ;
        RECT  14.25 7.15 15.10 8.90 ;
        RECT  14.25 8.00 15.15 8.90 ;
        RECT  14.60 2.60 15.30 4.30 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.40 19.35 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.85 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.40 6.30 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  8.55 5.40 9.55 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.40 5.40 2.55 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.15 2.50 11.00 ;
        RECT  4.65 9.15 5.35 11.00 ;
        RECT  9.00 7.20 9.70 11.00 ;
        RECT  12.90 7.20 13.60 11.00 ;
        RECT  15.60 7.20 16.30 11.00 ;
        RECT  18.45 7.75 19.15 11.00 ;
        RECT  18.05 10.10 20.55 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.40 ;
        RECT  8.85 2.00 9.55 4.35 ;
        RECT  11.55 2.00 12.25 4.35 ;
        RECT  13.25 2.00 13.95 4.30 ;
        RECT  15.95 2.00 16.65 4.30 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.30 7.15 8.20 7.50 ;
        RECT  0.45 3.70 0.95 9.85 ;
        RECT  0.45 3.70 1.15 4.40 ;
        RECT  0.45 8.15 1.15 9.85 ;
        RECT  0.45 7.00 2.85 7.50 ;
        RECT  2.15 7.00 2.85 7.70 ;
        RECT  3.30 3.70 3.80 9.85 ;
        RECT  3.30 8.20 4.00 9.85 ;
        RECT  4.30 7.00 5.00 7.70 ;
        RECT  5.15 2.65 5.85 4.20 ;
        RECT  3.30 3.70 5.85 4.20 ;
        RECT  3.30 8.20 6.50 8.70 ;
        RECT  6.00 8.20 6.50 9.85 ;
        RECT  6.00 9.15 6.70 9.85 ;
        RECT  7.15 2.45 7.85 3.15 ;
        RECT  5.15 2.65 7.85 3.15 ;
        RECT  7.50 3.65 8.00 8.85 ;
        RECT  4.30 7.00 8.00 7.50 ;
        RECT  7.50 3.65 8.20 4.35 ;
        RECT  7.50 7.15 8.20 8.85 ;
        RECT  10.20 3.70 10.90 4.40 ;
        RECT  10.40 3.70 10.90 5.30 ;
        RECT  11.55 4.80 12.05 10.55 ;
        RECT  11.35 7.15 12.05 10.55 ;
        RECT  10.40 4.80 14.05 5.30 ;
        RECT  13.35 4.80 14.05 5.50 ;
        RECT  17.10 7.70 17.60 10.55 ;
        RECT  17.30 3.80 17.60 10.55 ;
        RECT  16.90 9.85 17.60 10.55 ;
        RECT  17.30 3.80 17.80 8.40 ;
        RECT  17.10 7.70 17.80 8.40 ;
        RECT  17.30 6.75 20.50 7.25 ;
        RECT  19.45 3.60 20.15 4.30 ;
        RECT  17.30 3.80 20.15 4.30 ;
        RECT  19.80 6.75 20.50 8.40 ;
    END
END NA6I2X4
MACRO NA6I3X1
    CLASS CORE ;
    FOREIGN NA6I3X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.85 3.60 12.35 8.90 ;
        RECT  11.45 7.15 12.35 8.90 ;
        RECT  11.85 3.60 12.65 4.30 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 14.05 6.30 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.25 2.60 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.10 1.15 11.00 ;
        RECT  7.60 7.20 8.30 11.00 ;
        RECT  12.80 7.15 13.55 11.00 ;
        RECT  11.60 10.10 13.55 11.00 ;
        RECT  15.65 7.75 16.35 11.00 ;
        RECT  15.25 10.10 17.75 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.85 ;
        RECT  3.15 2.00 3.85 3.85 ;
        RECT  7.45 2.00 8.15 4.25 ;
        RECT  10.15 2.00 10.85 4.25 ;
        RECT  13.30 2.00 14.00 4.25 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.80 8.10 5.40 8.80 ;
        RECT  1.80 3.20 2.50 4.80 ;
        RECT  4.50 3.20 5.20 4.80 ;
        RECT  1.80 4.30 5.20 4.80 ;
        RECT  4.70 3.20 5.20 8.80 ;
        RECT  4.90 3.20 5.20 10.55 ;
        RECT  3.80 7.10 5.20 8.80 ;
        RECT  4.90 8.10 5.40 10.55 ;
        RECT  4.90 9.85 5.60 10.55 ;
        RECT  4.70 5.50 6.00 6.20 ;
        RECT  6.10 3.55 6.95 4.25 ;
        RECT  6.45 3.55 6.95 8.85 ;
        RECT  6.25 7.15 6.95 8.85 ;
        RECT  8.00 5.75 8.70 6.45 ;
        RECT  6.45 5.95 8.70 6.45 ;
        RECT  8.80 3.60 9.50 4.30 ;
        RECT  9.00 3.60 9.50 5.30 ;
        RECT  9.00 4.80 11.40 5.30 ;
        RECT  10.15 4.80 10.65 10.55 ;
        RECT  9.95 7.15 10.65 10.55 ;
        RECT  10.15 4.80 11.40 5.50 ;
        RECT  14.30 7.70 14.80 10.55 ;
        RECT  14.50 3.80 14.80 10.55 ;
        RECT  14.10 9.85 14.80 10.55 ;
        RECT  14.50 3.80 15.00 8.40 ;
        RECT  14.30 7.70 15.00 8.40 ;
        RECT  14.50 6.75 17.70 7.25 ;
        RECT  16.65 3.60 17.35 4.30 ;
        RECT  14.50 3.80 17.35 4.30 ;
        RECT  17.00 6.75 17.70 8.40 ;
    END
END NA6I3X1
MACRO NA6I3X2
    CLASS CORE ;
    FOREIGN NA6I3X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.80 2.70 12.15 10.55 ;
        RECT  11.45 7.15 12.15 10.55 ;
        RECT  11.80 2.70 12.30 9.20 ;
        RECT  11.45 7.15 12.30 9.20 ;
        RECT  11.45 8.00 12.35 9.20 ;
        RECT  11.80 2.70 12.50 4.30 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 14.05 6.30 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.25 2.60 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.10 1.15 11.00 ;
        RECT  7.60 7.20 8.30 11.00 ;
        RECT  12.80 7.20 13.55 11.00 ;
        RECT  15.65 7.75 16.35 11.00 ;
        RECT  15.25 10.10 17.75 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.85 ;
        RECT  3.15 2.00 3.85 3.85 ;
        RECT  7.45 2.00 8.15 4.25 ;
        RECT  10.15 2.00 10.85 4.25 ;
        RECT  13.15 2.00 13.85 4.25 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.80 8.10 5.40 8.80 ;
        RECT  1.80 3.20 2.50 4.80 ;
        RECT  4.50 3.20 5.20 4.80 ;
        RECT  1.80 4.30 5.20 4.80 ;
        RECT  4.70 3.20 5.20 8.80 ;
        RECT  4.90 3.20 5.20 10.55 ;
        RECT  3.80 7.10 5.20 8.80 ;
        RECT  4.90 8.10 5.40 10.55 ;
        RECT  4.90 9.85 5.60 10.55 ;
        RECT  4.70 5.50 6.00 6.20 ;
        RECT  6.10 3.55 6.95 4.25 ;
        RECT  6.45 3.55 6.95 8.85 ;
        RECT  6.25 7.15 6.95 8.85 ;
        RECT  8.00 5.75 8.70 6.45 ;
        RECT  6.45 5.95 8.70 6.45 ;
        RECT  8.80 3.60 9.50 4.30 ;
        RECT  9.00 3.60 9.50 5.30 ;
        RECT  9.00 4.80 11.35 5.30 ;
        RECT  10.15 4.80 10.65 10.55 ;
        RECT  9.95 7.15 10.65 10.55 ;
        RECT  10.15 4.80 11.35 5.50 ;
        RECT  14.30 7.70 14.80 10.55 ;
        RECT  14.50 3.80 14.80 10.55 ;
        RECT  14.10 9.85 14.80 10.55 ;
        RECT  14.50 3.80 15.00 8.40 ;
        RECT  14.30 7.70 15.00 8.40 ;
        RECT  14.50 6.75 17.70 7.25 ;
        RECT  16.65 3.60 17.35 4.30 ;
        RECT  14.50 3.80 17.35 4.30 ;
        RECT  17.00 6.75 17.70 8.40 ;
    END
END NA6I3X2
MACRO NA6I3X4
    CLASS CORE ;
    FOREIGN NA6I3X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  13.20 2.70 13.55 10.55 ;
        RECT  12.85 7.15 13.55 10.55 ;
        RECT  13.20 2.70 13.70 9.20 ;
        RECT  12.85 7.15 13.70 9.20 ;
        RECT  12.85 8.00 13.75 9.20 ;
        RECT  13.20 2.70 13.90 4.30 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.40 19.35 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.45 6.30 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.25 2.60 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.10 1.15 11.00 ;
        RECT  7.60 7.20 8.30 11.00 ;
        RECT  11.50 7.20 12.20 11.00 ;
        RECT  14.20 7.20 14.90 11.00 ;
        RECT  17.05 7.75 17.75 11.00 ;
        RECT  16.65 10.10 19.15 11.00 ;
        RECT  0.00 11.00 19.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.85 ;
        RECT  3.15 2.00 3.85 3.85 ;
        RECT  7.45 2.00 8.15 4.25 ;
        RECT  10.15 2.00 10.85 4.25 ;
        RECT  11.85 2.00 12.55 4.25 ;
        RECT  14.55 2.00 15.25 4.25 ;
        RECT  0.00 0.00 19.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.80 8.10 5.40 8.80 ;
        RECT  1.80 3.20 2.50 4.80 ;
        RECT  4.50 3.20 5.20 4.80 ;
        RECT  1.80 4.30 5.20 4.80 ;
        RECT  4.70 3.20 5.20 8.80 ;
        RECT  4.90 3.20 5.20 10.55 ;
        RECT  3.80 7.10 5.20 8.80 ;
        RECT  4.90 8.10 5.40 10.55 ;
        RECT  4.90 9.85 5.60 10.55 ;
        RECT  4.70 5.50 6.00 6.20 ;
        RECT  6.10 3.55 6.95 4.25 ;
        RECT  6.45 3.55 6.95 8.85 ;
        RECT  6.25 7.15 6.95 8.85 ;
        RECT  8.00 5.75 8.70 6.45 ;
        RECT  6.45 5.95 8.70 6.45 ;
        RECT  8.80 3.60 9.50 4.30 ;
        RECT  9.00 3.60 9.50 5.30 ;
        RECT  10.15 4.80 10.65 10.55 ;
        RECT  9.95 7.15 10.65 10.55 ;
        RECT  9.00 4.80 12.65 5.30 ;
        RECT  11.95 4.80 12.65 5.50 ;
        RECT  15.70 7.70 16.20 10.55 ;
        RECT  15.90 3.80 16.20 10.55 ;
        RECT  15.50 9.85 16.20 10.55 ;
        RECT  15.90 3.80 16.40 8.40 ;
        RECT  15.70 7.70 16.40 8.40 ;
        RECT  15.90 6.75 19.10 7.25 ;
        RECT  18.05 3.60 18.75 4.30 ;
        RECT  15.90 3.80 18.75 4.30 ;
        RECT  18.40 6.75 19.10 8.40 ;
    END
END NA6I3X4
MACRO NA6I4X1
    CLASS CORE ;
    FOREIGN NA6I4X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.85 3.60 12.35 8.90 ;
        RECT  11.45 7.15 12.35 8.90 ;
        RECT  11.85 3.60 12.65 4.30 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END E
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END DN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.25 2.60 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.10 1.15 11.00 ;
        RECT  7.60 7.20 8.30 11.00 ;
        RECT  12.80 7.15 13.55 11.00 ;
        RECT  11.60 10.10 13.55 11.00 ;
        RECT  15.65 7.75 16.35 11.00 ;
        RECT  19.85 7.15 20.55 11.00 ;
        RECT  15.25 10.10 20.55 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.85 ;
        RECT  3.15 2.00 3.85 3.85 ;
        RECT  7.45 2.00 8.15 4.25 ;
        RECT  10.15 2.00 10.85 4.25 ;
        RECT  13.30 2.00 14.00 4.25 ;
        RECT  19.85 2.00 20.55 4.30 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.80 8.10 5.40 8.80 ;
        RECT  1.80 3.20 2.50 4.80 ;
        RECT  4.50 3.20 5.20 4.80 ;
        RECT  1.80 4.30 5.20 4.80 ;
        RECT  4.70 3.20 5.20 8.80 ;
        RECT  4.90 3.20 5.20 10.55 ;
        RECT  3.80 7.10 5.20 8.80 ;
        RECT  4.90 8.10 5.40 10.55 ;
        RECT  4.90 9.85 5.60 10.55 ;
        RECT  4.70 5.50 6.00 6.20 ;
        RECT  6.10 3.55 6.95 4.25 ;
        RECT  6.45 3.55 6.95 8.85 ;
        RECT  6.25 7.15 6.95 8.85 ;
        RECT  8.00 5.75 8.70 6.45 ;
        RECT  6.45 5.95 8.70 6.45 ;
        RECT  8.80 3.60 9.50 4.30 ;
        RECT  9.00 3.60 9.50 5.30 ;
        RECT  9.00 4.80 11.40 5.30 ;
        RECT  10.15 4.80 10.65 10.55 ;
        RECT  9.95 7.15 10.65 10.55 ;
        RECT  10.15 4.80 11.40 5.50 ;
        RECT  14.30 7.70 14.80 10.55 ;
        RECT  14.50 3.80 14.80 10.55 ;
        RECT  14.10 9.85 14.80 10.55 ;
        RECT  14.50 3.80 15.00 8.40 ;
        RECT  14.30 7.70 15.00 8.40 ;
        RECT  14.50 6.75 17.70 7.25 ;
        RECT  16.65 3.60 17.35 4.30 ;
        RECT  14.50 3.80 17.35 4.30 ;
        RECT  17.00 6.75 17.70 8.40 ;
        RECT  18.15 2.45 19.00 3.15 ;
        RECT  18.50 2.45 19.00 8.85 ;
        RECT  18.50 3.60 19.20 4.30 ;
        RECT  18.50 7.15 19.20 8.85 ;
    END
END NA6I4X1
MACRO NA6I4X2
    CLASS CORE ;
    FOREIGN NA6I4X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.80 2.70 12.15 10.55 ;
        RECT  11.45 7.15 12.15 10.55 ;
        RECT  11.80 2.70 12.30 9.20 ;
        RECT  11.45 7.15 12.30 9.20 ;
        RECT  11.45 8.00 12.35 9.20 ;
        RECT  11.80 2.70 12.50 4.30 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END E
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END DN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.25 2.60 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.10 1.15 11.00 ;
        RECT  7.60 7.20 8.30 11.00 ;
        RECT  12.80 7.15 13.50 11.00 ;
        RECT  15.65 7.75 16.35 11.00 ;
        RECT  19.85 7.15 20.55 11.00 ;
        RECT  15.25 10.10 20.55 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.85 ;
        RECT  3.15 2.00 3.85 3.85 ;
        RECT  7.45 2.00 8.15 4.25 ;
        RECT  10.15 2.00 10.85 4.25 ;
        RECT  13.15 2.00 13.85 4.25 ;
        RECT  19.85 2.00 20.55 4.30 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.80 8.10 5.40 8.80 ;
        RECT  1.80 3.20 2.50 4.80 ;
        RECT  4.50 3.20 5.20 4.80 ;
        RECT  1.80 4.30 5.20 4.80 ;
        RECT  4.70 3.20 5.20 8.80 ;
        RECT  4.90 3.20 5.20 10.55 ;
        RECT  3.80 7.10 5.20 8.80 ;
        RECT  4.90 8.10 5.40 10.55 ;
        RECT  4.90 9.85 5.60 10.55 ;
        RECT  4.70 5.50 6.00 6.20 ;
        RECT  6.10 3.55 6.95 4.25 ;
        RECT  6.45 3.55 6.95 8.85 ;
        RECT  6.25 7.15 6.95 8.85 ;
        RECT  8.00 5.75 8.70 6.45 ;
        RECT  6.45 5.95 8.70 6.45 ;
        RECT  8.80 3.60 9.50 4.30 ;
        RECT  9.00 3.60 9.50 5.30 ;
        RECT  9.00 4.80 11.35 5.30 ;
        RECT  10.15 4.80 10.65 10.55 ;
        RECT  9.95 7.15 10.65 10.55 ;
        RECT  10.15 4.80 11.35 5.50 ;
        RECT  14.30 7.70 14.80 10.55 ;
        RECT  14.50 3.80 14.80 10.55 ;
        RECT  14.10 9.85 14.80 10.55 ;
        RECT  14.50 3.80 15.00 8.40 ;
        RECT  14.30 7.70 15.00 8.40 ;
        RECT  14.50 6.75 17.70 7.25 ;
        RECT  16.65 3.60 17.35 4.30 ;
        RECT  14.50 3.80 17.35 4.30 ;
        RECT  17.00 6.75 17.70 8.40 ;
        RECT  18.15 2.45 19.00 3.15 ;
        RECT  18.50 2.45 19.00 8.85 ;
        RECT  18.50 3.60 19.20 4.30 ;
        RECT  18.50 7.15 19.20 8.85 ;
    END
END NA6I4X2
MACRO NA6I4X4
    CLASS CORE ;
    FOREIGN NA6I4X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  13.20 2.70 13.55 10.55 ;
        RECT  12.85 7.15 13.55 10.55 ;
        RECT  13.20 2.70 13.70 9.20 ;
        RECT  12.85 7.15 13.70 9.20 ;
        RECT  12.85 8.00 13.75 9.20 ;
        RECT  13.20 2.70 13.90 4.30 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.40 19.35 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END E
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  21.25 5.40 22.15 6.30 ;
        END
    END DN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.25 2.60 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.10 1.15 11.00 ;
        RECT  7.60 7.20 8.30 11.00 ;
        RECT  11.50 7.15 12.20 11.00 ;
        RECT  14.20 7.15 14.90 11.00 ;
        RECT  17.05 7.75 17.75 11.00 ;
        RECT  21.25 7.15 21.95 11.00 ;
        RECT  16.65 10.10 21.95 11.00 ;
        RECT  0.00 11.00 22.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.85 ;
        RECT  3.15 2.00 3.85 3.85 ;
        RECT  7.45 2.00 8.15 4.25 ;
        RECT  10.15 2.00 10.85 4.25 ;
        RECT  11.85 2.00 12.55 4.25 ;
        RECT  14.55 2.00 15.25 4.25 ;
        RECT  21.25 2.00 21.95 4.30 ;
        RECT  0.00 0.00 22.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.80 8.10 5.40 8.80 ;
        RECT  1.80 3.20 2.50 4.80 ;
        RECT  4.50 3.20 5.20 4.80 ;
        RECT  1.80 4.30 5.20 4.80 ;
        RECT  4.70 3.20 5.20 8.80 ;
        RECT  4.90 3.20 5.20 10.55 ;
        RECT  3.80 7.10 5.20 8.80 ;
        RECT  4.90 8.10 5.40 10.55 ;
        RECT  4.90 9.85 5.60 10.55 ;
        RECT  4.70 5.50 6.00 6.20 ;
        RECT  6.10 3.55 6.95 4.25 ;
        RECT  6.45 3.55 6.95 8.85 ;
        RECT  6.25 7.15 6.95 8.85 ;
        RECT  8.00 5.75 8.70 6.45 ;
        RECT  6.45 5.95 8.70 6.45 ;
        RECT  8.80 3.60 9.50 4.30 ;
        RECT  9.00 3.60 9.50 5.30 ;
        RECT  10.15 4.80 10.65 10.55 ;
        RECT  9.95 7.15 10.65 10.55 ;
        RECT  9.00 4.80 12.65 5.30 ;
        RECT  11.95 4.80 12.65 5.50 ;
        RECT  15.70 7.70 16.20 10.55 ;
        RECT  15.90 3.80 16.20 10.55 ;
        RECT  15.50 9.85 16.20 10.55 ;
        RECT  15.90 3.80 16.40 8.40 ;
        RECT  15.70 7.70 16.40 8.40 ;
        RECT  15.90 6.75 19.10 7.25 ;
        RECT  18.05 3.60 18.75 4.30 ;
        RECT  15.90 3.80 18.75 4.30 ;
        RECT  18.40 6.75 19.10 8.40 ;
        RECT  19.55 2.45 20.40 3.15 ;
        RECT  19.90 2.45 20.40 8.85 ;
        RECT  19.90 3.60 20.60 4.30 ;
        RECT  19.90 7.15 20.60 8.85 ;
    END
END NA6I4X4
MACRO NA6I5X1
    CLASS CORE ;
    FOREIGN NA6I5X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.85 3.60 12.35 8.90 ;
        RECT  11.45 7.15 12.35 8.90 ;
        RECT  11.85 3.60 12.65 4.30 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END F
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  18.45 9.30 19.35 10.20 ;
        END
    END EN
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END DN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.25 2.60 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.10 1.15 11.00 ;
        RECT  7.60 7.20 8.30 11.00 ;
        RECT  12.80 7.15 13.55 11.00 ;
        RECT  11.60 10.10 13.55 11.00 ;
        RECT  15.65 7.75 16.35 11.00 ;
        RECT  15.50 10.10 18.00 11.00 ;
        RECT  19.85 7.25 20.55 11.00 ;
        RECT  19.85 10.10 21.95 11.00 ;
        RECT  0.00 11.00 22.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.85 ;
        RECT  3.15 2.00 3.85 3.85 ;
        RECT  7.45 2.00 8.15 4.25 ;
        RECT  10.15 2.00 10.85 4.25 ;
        RECT  13.30 2.00 14.00 4.25 ;
        RECT  19.60 2.00 20.30 4.30 ;
        RECT  0.00 0.00 22.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.80 8.10 5.40 8.80 ;
        RECT  1.80 3.20 2.50 4.80 ;
        RECT  4.50 3.20 5.20 4.80 ;
        RECT  1.80 4.30 5.20 4.80 ;
        RECT  4.70 3.20 5.20 8.80 ;
        RECT  4.90 3.20 5.20 10.55 ;
        RECT  3.80 7.10 5.20 8.80 ;
        RECT  4.90 8.10 5.40 10.55 ;
        RECT  4.90 9.85 5.60 10.55 ;
        RECT  4.70 5.50 6.00 6.20 ;
        RECT  6.10 3.55 6.95 4.25 ;
        RECT  6.45 3.55 6.95 8.85 ;
        RECT  6.25 7.15 6.95 8.85 ;
        RECT  8.00 5.75 8.70 6.45 ;
        RECT  6.45 5.95 8.70 6.45 ;
        RECT  8.80 3.60 9.50 4.30 ;
        RECT  9.00 3.60 9.50 5.30 ;
        RECT  9.00 4.80 11.40 5.30 ;
        RECT  10.15 4.80 10.65 10.55 ;
        RECT  9.95 7.15 10.65 10.55 ;
        RECT  10.15 4.80 11.40 5.50 ;
        RECT  14.30 7.70 14.80 10.55 ;
        RECT  14.50 3.50 14.80 10.55 ;
        RECT  14.10 9.85 14.80 10.55 ;
        RECT  14.50 3.50 15.00 8.40 ;
        RECT  14.30 7.70 15.00 8.40 ;
        RECT  15.65 4.45 16.15 6.25 ;
        RECT  15.45 5.55 16.15 6.25 ;
        RECT  14.50 6.75 17.70 7.25 ;
        RECT  16.65 3.30 17.35 4.00 ;
        RECT  14.50 3.50 17.35 4.00 ;
        RECT  17.00 6.75 17.70 8.40 ;
        RECT  18.25 3.60 19.00 4.95 ;
        RECT  15.65 4.45 19.00 4.95 ;
        RECT  18.50 3.60 19.00 8.85 ;
        RECT  18.50 7.25 19.20 8.85 ;
        RECT  20.95 3.60 21.70 4.30 ;
        RECT  21.20 2.45 21.70 8.85 ;
        RECT  21.20 7.25 21.90 8.85 ;
        RECT  21.20 2.45 22.00 3.15 ;
    END
END NA6I5X1
MACRO NA6I5X2
    CLASS CORE ;
    FOREIGN NA6I5X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.80 2.70 12.15 10.55 ;
        RECT  11.45 7.15 12.15 10.55 ;
        RECT  11.80 2.70 12.30 9.20 ;
        RECT  11.45 7.15 12.30 9.20 ;
        RECT  11.45 8.00 12.35 9.20 ;
        RECT  11.80 2.70 12.50 4.30 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END F
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  18.45 9.30 19.35 10.20 ;
        END
    END EN
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END DN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.25 2.60 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.10 1.15 11.00 ;
        RECT  7.60 7.20 8.30 11.00 ;
        RECT  12.80 7.15 13.50 11.00 ;
        RECT  15.65 7.75 16.35 11.00 ;
        RECT  15.50 10.10 18.00 11.00 ;
        RECT  19.85 7.25 20.55 11.00 ;
        RECT  19.85 10.10 21.95 11.00 ;
        RECT  0.00 11.00 22.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.85 ;
        RECT  3.15 2.00 3.85 3.85 ;
        RECT  7.45 2.00 8.15 4.25 ;
        RECT  10.15 2.00 10.85 4.25 ;
        RECT  13.15 2.00 13.85 4.25 ;
        RECT  19.60 2.00 20.30 4.30 ;
        RECT  0.00 0.00 22.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.80 8.10 5.40 8.80 ;
        RECT  1.80 3.20 2.50 4.80 ;
        RECT  4.50 3.20 5.20 4.80 ;
        RECT  1.80 4.30 5.20 4.80 ;
        RECT  4.70 3.20 5.20 8.80 ;
        RECT  4.90 3.20 5.20 10.55 ;
        RECT  3.80 7.10 5.20 8.80 ;
        RECT  4.90 8.10 5.40 10.55 ;
        RECT  4.90 9.85 5.60 10.55 ;
        RECT  4.70 5.50 6.00 6.20 ;
        RECT  6.10 3.55 6.95 4.25 ;
        RECT  6.45 3.55 6.95 8.85 ;
        RECT  6.25 7.15 6.95 8.85 ;
        RECT  8.00 5.75 8.70 6.45 ;
        RECT  6.45 5.95 8.70 6.45 ;
        RECT  8.80 3.60 9.50 4.30 ;
        RECT  9.00 3.60 9.50 5.30 ;
        RECT  9.00 4.80 11.35 5.30 ;
        RECT  10.15 4.80 10.65 10.55 ;
        RECT  9.95 7.15 10.65 10.55 ;
        RECT  10.15 4.80 11.35 5.50 ;
        RECT  14.30 7.70 14.80 10.55 ;
        RECT  14.50 3.50 14.80 10.55 ;
        RECT  14.10 9.85 14.80 10.55 ;
        RECT  14.50 3.50 15.00 8.40 ;
        RECT  14.30 7.70 15.00 8.40 ;
        RECT  15.65 4.45 16.15 6.25 ;
        RECT  15.45 5.55 16.15 6.25 ;
        RECT  14.50 6.75 17.70 7.25 ;
        RECT  16.65 3.30 17.35 4.00 ;
        RECT  14.50 3.50 17.35 4.00 ;
        RECT  17.00 6.75 17.70 8.40 ;
        RECT  18.25 3.60 19.00 4.95 ;
        RECT  15.65 4.45 19.00 4.95 ;
        RECT  18.50 3.60 19.00 8.85 ;
        RECT  18.50 7.25 19.20 8.85 ;
        RECT  20.95 3.60 21.70 4.30 ;
        RECT  21.20 2.45 21.70 8.85 ;
        RECT  21.20 7.25 21.90 8.85 ;
        RECT  21.20 2.45 22.00 3.15 ;
    END
END NA6I5X2
MACRO NA6I5X4
    CLASS CORE ;
    FOREIGN NA6I5X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  13.20 2.70 13.55 10.55 ;
        RECT  12.85 7.15 13.55 10.55 ;
        RECT  13.20 2.70 13.70 9.20 ;
        RECT  12.85 7.15 13.70 9.20 ;
        RECT  12.85 8.00 13.75 9.20 ;
        RECT  13.20 2.70 13.90 4.30 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.40 19.35 6.30 ;
        END
    END F
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  19.85 9.30 20.75 10.20 ;
        END
    END EN
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  21.25 5.40 22.15 6.30 ;
        END
    END DN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.25 2.60 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.10 1.15 11.00 ;
        RECT  7.60 7.20 8.30 11.00 ;
        RECT  11.50 7.15 12.20 11.00 ;
        RECT  14.20 7.15 14.90 11.00 ;
        RECT  17.05 7.75 17.75 11.00 ;
        RECT  16.90 10.10 19.40 11.00 ;
        RECT  21.25 7.25 21.95 11.00 ;
        RECT  21.25 10.10 23.35 11.00 ;
        RECT  0.00 11.00 23.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.85 ;
        RECT  3.15 2.00 3.85 3.85 ;
        RECT  7.45 2.00 8.15 4.25 ;
        RECT  10.15 2.00 10.85 4.25 ;
        RECT  11.85 2.00 12.55 4.25 ;
        RECT  14.55 2.00 15.25 4.25 ;
        RECT  21.00 2.00 21.70 4.30 ;
        RECT  0.00 0.00 23.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.80 8.10 5.40 8.80 ;
        RECT  1.80 3.20 2.50 4.80 ;
        RECT  4.50 3.20 5.20 4.80 ;
        RECT  1.80 4.30 5.20 4.80 ;
        RECT  4.70 3.20 5.20 8.80 ;
        RECT  4.90 3.20 5.20 10.55 ;
        RECT  3.80 7.10 5.20 8.80 ;
        RECT  4.90 8.10 5.40 10.55 ;
        RECT  4.90 9.85 5.60 10.55 ;
        RECT  4.70 5.50 6.00 6.20 ;
        RECT  6.10 3.55 6.95 4.25 ;
        RECT  6.45 3.55 6.95 8.85 ;
        RECT  6.25 7.15 6.95 8.85 ;
        RECT  8.00 5.75 8.70 6.45 ;
        RECT  6.45 5.95 8.70 6.45 ;
        RECT  8.80 3.60 9.50 4.30 ;
        RECT  9.00 3.60 9.50 5.30 ;
        RECT  10.15 4.80 10.65 10.55 ;
        RECT  9.95 7.15 10.65 10.55 ;
        RECT  9.00 4.80 12.65 5.30 ;
        RECT  11.95 4.80 12.65 5.50 ;
        RECT  15.70 7.70 16.20 10.55 ;
        RECT  15.90 3.50 16.20 10.55 ;
        RECT  15.50 9.85 16.20 10.55 ;
        RECT  15.90 3.50 16.40 8.40 ;
        RECT  15.70 7.70 16.40 8.40 ;
        RECT  17.05 4.45 17.55 6.25 ;
        RECT  16.85 5.55 17.55 6.25 ;
        RECT  15.90 6.75 19.10 7.25 ;
        RECT  18.05 3.30 18.75 4.00 ;
        RECT  15.90 3.50 18.75 4.00 ;
        RECT  18.40 6.75 19.10 8.40 ;
        RECT  19.65 3.60 20.40 4.95 ;
        RECT  17.05 4.45 20.40 4.95 ;
        RECT  19.90 3.60 20.40 8.85 ;
        RECT  19.90 7.25 20.60 8.85 ;
        RECT  22.35 3.60 23.10 4.30 ;
        RECT  22.60 2.45 23.10 8.85 ;
        RECT  22.60 7.25 23.30 8.85 ;
        RECT  22.60 2.45 23.40 3.15 ;
    END
END NA6I5X4
MACRO NA6X1
    CLASS CORE ;
    FOREIGN NA6X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  9.05 3.60 9.55 9.20 ;
        RECT  8.65 7.10 9.55 9.20 ;
        RECT  9.05 3.60 9.85 4.30 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 11.25 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  0.25 6.70 1.15 7.60 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.55 7.60 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 4.45 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 9.15 2.55 11.00 ;
        RECT  4.70 7.20 5.40 11.00 ;
        RECT  10.00 7.45 10.75 11.00 ;
        RECT  9.15 10.10 10.75 11.00 ;
        RECT  12.85 8.15 13.55 11.00 ;
        RECT  12.85 10.10 14.90 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  4.20 2.00 4.90 3.65 ;
        RECT  6.90 2.00 7.60 3.65 ;
        RECT  10.50 2.00 11.20 4.25 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.85 2.80 1.55 3.50 ;
        RECT  0.50 8.20 1.20 9.85 ;
        RECT  1.05 2.80 1.55 6.05 ;
        RECT  0.50 8.20 3.90 8.70 ;
        RECT  3.40 5.55 3.90 9.85 ;
        RECT  3.20 8.20 3.90 9.85 ;
        RECT  1.05 5.55 5.85 6.05 ;
        RECT  5.55 3.00 6.25 3.70 ;
        RECT  5.15 5.55 5.85 6.25 ;
        RECT  5.75 3.00 6.25 4.75 ;
        RECT  5.75 4.25 8.35 4.75 ;
        RECT  7.25 4.25 7.75 10.55 ;
        RECT  7.05 7.15 7.75 10.55 ;
        RECT  7.25 4.25 8.35 4.95 ;
        RECT  11.70 3.80 12.20 10.55 ;
        RECT  11.50 8.10 12.20 10.55 ;
        RECT  11.70 7.15 14.90 7.65 ;
        RECT  13.85 3.60 14.55 4.30 ;
        RECT  11.70 3.80 14.55 4.30 ;
        RECT  14.20 7.15 14.90 8.80 ;
    END
END NA6X1
MACRO NA6X2
    CLASS CORE ;
    FOREIGN NA6X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.65 2.60 9.15 10.55 ;
        RECT  8.65 2.60 9.35 4.35 ;
        RECT  8.65 7.15 9.35 10.55 ;
        RECT  8.65 8.00 9.55 8.90 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 11.25 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  0.25 6.70 1.15 7.60 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.55 7.60 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 4.45 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 9.05 2.55 11.00 ;
        RECT  4.70 7.20 5.40 11.00 ;
        RECT  10.00 7.15 10.70 11.00 ;
        RECT  12.85 7.70 13.55 11.00 ;
        RECT  11.50 10.10 14.95 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  4.20 2.00 4.90 3.65 ;
        RECT  6.90 2.00 7.60 3.65 ;
        RECT  10.00 2.00 10.70 4.35 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.85 2.80 1.55 3.50 ;
        RECT  0.70 8.10 1.20 9.75 ;
        RECT  0.50 9.05 1.20 9.75 ;
        RECT  1.05 2.80 1.55 6.05 ;
        RECT  0.70 8.10 3.70 8.60 ;
        RECT  3.20 5.55 3.70 9.75 ;
        RECT  3.20 9.05 3.90 9.75 ;
        RECT  1.05 5.55 5.85 6.05 ;
        RECT  5.55 3.00 6.25 3.70 ;
        RECT  5.15 5.55 5.85 6.25 ;
        RECT  5.75 3.00 6.25 5.00 ;
        RECT  5.75 4.50 8.20 5.00 ;
        RECT  7.25 4.50 7.75 10.55 ;
        RECT  7.05 7.15 7.75 10.55 ;
        RECT  7.25 4.50 8.20 5.20 ;
        RECT  11.70 3.80 12.20 8.40 ;
        RECT  11.50 7.70 12.20 8.40 ;
        RECT  13.50 3.60 14.45 4.30 ;
        RECT  11.70 6.75 14.70 7.25 ;
        RECT  13.95 2.45 14.45 4.30 ;
        RECT  11.70 3.80 14.45 4.30 ;
        RECT  14.20 6.75 14.70 8.40 ;
        RECT  13.95 2.45 14.90 3.15 ;
        RECT  14.20 7.70 14.90 8.40 ;
    END
END NA6X2
MACRO NA6X3
    CLASS CORE ;
    FOREIGN NA6X3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.75 2.45 9.25 10.55 ;
        RECT  8.55 7.15 9.25 10.55 ;
        RECT  8.65 2.45 9.35 4.35 ;
        RECT  8.55 9.30 9.55 10.55 ;
        RECT  8.55 9.85 10.20 10.55 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 11.25 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  0.25 6.70 1.15 7.60 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.55 7.60 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 4.45 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 9.00 2.55 11.00 ;
        RECT  4.70 7.20 5.40 11.00 ;
        RECT  9.90 7.15 10.60 9.00 ;
        RECT  9.90 8.50 11.55 9.00 ;
        RECT  10.85 8.50 11.55 11.00 ;
        RECT  12.90 7.70 13.60 11.00 ;
        RECT  12.45 10.10 14.95 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  4.20 2.00 4.90 3.65 ;
        RECT  6.90 2.00 7.60 3.65 ;
        RECT  10.00 2.00 10.70 4.35 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.85 3.05 1.55 3.75 ;
        RECT  0.70 8.05 1.20 9.70 ;
        RECT  0.50 9.00 1.20 9.70 ;
        RECT  1.05 3.05 1.55 6.05 ;
        RECT  0.70 8.05 3.70 8.55 ;
        RECT  3.20 5.55 3.70 9.70 ;
        RECT  3.20 9.00 3.90 9.70 ;
        RECT  1.05 5.55 5.85 6.05 ;
        RECT  5.55 3.00 6.25 3.70 ;
        RECT  5.15 5.55 5.85 6.25 ;
        RECT  5.75 3.00 6.25 5.00 ;
        RECT  5.75 4.50 8.20 5.00 ;
        RECT  7.25 4.50 7.75 10.55 ;
        RECT  7.05 7.15 7.75 10.55 ;
        RECT  7.25 4.50 8.20 5.20 ;
        RECT  11.70 3.80 12.20 7.85 ;
        RECT  11.40 7.15 12.20 7.85 ;
        RECT  13.50 3.60 14.70 4.30 ;
        RECT  11.70 6.75 14.75 7.25 ;
        RECT  11.40 7.15 14.75 7.25 ;
        RECT  14.20 2.45 14.70 4.30 ;
        RECT  11.70 3.80 14.70 4.30 ;
        RECT  14.25 6.75 14.75 8.40 ;
        RECT  14.20 2.45 14.90 3.15 ;
        RECT  14.25 7.70 14.95 8.40 ;
    END
END NA6X3
MACRO NA6X4
    CLASS CORE ;
    FOREIGN NA6X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.75 4.10 9.25 10.55 ;
        RECT  8.80 2.55 9.25 10.55 ;
        RECT  8.55 7.15 9.25 10.55 ;
        RECT  8.80 2.55 9.55 5.00 ;
        RECT  8.65 4.10 9.55 5.00 ;
        RECT  8.55 9.85 11.10 10.55 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 11.25 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  0.25 6.70 1.15 7.60 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.55 7.60 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 4.25 7.60 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 9.00 2.55 11.00 ;
        RECT  4.70 9.00 5.40 11.00 ;
        RECT  9.90 7.20 10.60 9.20 ;
        RECT  11.75 8.60 12.45 11.00 ;
        RECT  12.90 7.70 13.60 9.20 ;
        RECT  9.90 8.60 13.60 9.20 ;
        RECT  13.35 10.10 14.95 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  4.20 2.00 4.90 4.40 ;
        RECT  6.90 2.00 7.60 4.40 ;
        RECT  10.15 2.00 10.85 4.50 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.85 3.50 1.55 4.20 ;
        RECT  0.70 8.05 1.20 9.60 ;
        RECT  0.50 8.90 1.20 9.60 ;
        RECT  1.05 3.50 1.55 5.65 ;
        RECT  3.20 8.05 3.90 9.60 ;
        RECT  1.05 5.15 5.20 5.65 ;
        RECT  4.70 5.15 5.20 8.55 ;
        RECT  0.70 8.05 5.20 8.55 ;
        RECT  5.55 3.75 6.25 4.45 ;
        RECT  4.70 5.80 5.80 6.50 ;
        RECT  5.75 3.75 6.25 5.35 ;
        RECT  5.75 4.85 8.20 5.35 ;
        RECT  7.25 4.85 7.75 10.55 ;
        RECT  7.05 8.05 7.75 10.55 ;
        RECT  7.25 4.85 8.20 5.55 ;
        RECT  11.70 3.80 12.20 7.90 ;
        RECT  11.40 7.20 12.20 7.90 ;
        RECT  13.65 3.60 14.50 4.30 ;
        RECT  11.70 6.75 14.75 7.25 ;
        RECT  11.40 7.20 14.75 7.25 ;
        RECT  14.00 2.45 14.50 4.30 ;
        RECT  11.70 3.80 14.50 4.30 ;
        RECT  14.25 6.75 14.75 8.40 ;
        RECT  14.25 7.70 14.95 8.40 ;
        RECT  14.00 2.45 15.05 3.15 ;
    END
END NA6X4
MACRO NA7X1
    CLASS CORE ;
    FOREIGN NA7X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  9.55 3.80 10.95 4.50 ;
        RECT  10.05 3.80 10.55 8.95 ;
        RECT  10.05 7.35 10.80 8.95 ;
        RECT  10.05 3.80 10.95 5.00 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  14.10 5.40 15.15 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  12.85 9.30 13.75 10.20 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  15.65 9.30 16.55 10.20 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.70 2.50 11.00 ;
        RECT  0.45 10.10 3.85 11.00 ;
        RECT  4.65 7.70 5.35 11.00 ;
        RECT  11.40 7.35 12.10 11.00 ;
        RECT  9.85 10.10 12.10 11.00 ;
        RECT  14.25 7.35 14.95 11.00 ;
        RECT  16.95 7.35 17.75 8.05 ;
        RECT  17.05 7.35 17.75 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.80 2.00 4.50 3.85 ;
        RECT  6.50 2.00 7.20 3.85 ;
        RECT  9.55 2.00 10.25 3.15 ;
        RECT  14.45 2.00 15.15 4.45 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 6.75 1.15 8.40 ;
        RECT  0.45 2.95 2.25 3.65 ;
        RECT  1.75 2.95 2.25 4.95 ;
        RECT  3.15 6.75 3.85 8.40 ;
        RECT  1.75 4.45 4.90 4.95 ;
        RECT  4.40 4.45 4.90 7.25 ;
        RECT  0.45 6.75 4.90 7.25 ;
        RECT  5.15 3.15 5.85 3.85 ;
        RECT  4.40 5.50 5.80 6.20 ;
        RECT  5.35 3.15 5.85 4.95 ;
        RECT  7.85 3.15 8.55 4.95 ;
        RECT  8.00 3.15 8.55 10.55 ;
        RECT  5.35 4.45 8.55 4.95 ;
        RECT  8.00 4.95 8.70 10.55 ;
        RECT  8.00 4.95 9.10 5.65 ;
        RECT  11.30 2.45 12.60 3.15 ;
        RECT  12.10 2.45 12.60 4.45 ;
        RECT  12.10 3.75 13.40 4.45 ;
        RECT  12.90 3.75 13.40 8.05 ;
        RECT  12.90 7.35 13.60 8.05 ;
        RECT  15.80 3.95 16.30 8.05 ;
        RECT  15.60 7.35 16.30 8.05 ;
        RECT  16.80 2.45 17.50 4.45 ;
        RECT  15.80 3.95 17.50 4.45 ;
        RECT  16.80 2.45 17.85 3.15 ;
    END
END NA7X1
MACRO NA7X2
    CLASS CORE ;
    FOREIGN NA7X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.05 3.80 10.55 10.55 ;
        RECT  10.05 7.15 10.80 10.55 ;
        RECT  10.05 8.00 10.95 8.90 ;
        RECT  9.70 3.80 11.30 4.50 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  14.10 5.25 15.15 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.45 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  15.65 9.30 16.55 10.20 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.70 2.50 11.00 ;
        RECT  0.45 10.10 3.85 11.00 ;
        RECT  4.65 7.70 5.35 11.00 ;
        RECT  11.40 7.35 12.10 11.00 ;
        RECT  14.25 7.15 14.95 11.00 ;
        RECT  16.95 7.15 17.75 7.85 ;
        RECT  17.05 7.15 17.75 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.80 2.00 4.50 3.85 ;
        RECT  6.50 2.00 7.20 3.85 ;
        RECT  9.65 2.00 11.25 3.15 ;
        RECT  14.50 2.00 15.20 4.45 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 6.75 1.15 8.40 ;
        RECT  0.45 2.95 2.25 3.65 ;
        RECT  1.75 2.95 2.25 4.95 ;
        RECT  3.15 6.75 3.85 8.40 ;
        RECT  1.75 4.45 4.90 4.95 ;
        RECT  4.40 4.45 4.90 7.25 ;
        RECT  0.45 6.75 4.90 7.25 ;
        RECT  5.15 3.15 5.85 3.85 ;
        RECT  4.40 5.50 5.80 6.20 ;
        RECT  5.35 3.15 5.85 4.95 ;
        RECT  7.85 3.15 8.55 4.95 ;
        RECT  8.00 3.15 8.55 10.55 ;
        RECT  5.35 4.45 8.55 4.95 ;
        RECT  8.00 4.95 8.70 10.55 ;
        RECT  8.00 4.95 9.10 5.65 ;
        RECT  12.15 3.75 13.40 4.45 ;
        RECT  12.90 3.75 13.40 10.55 ;
        RECT  12.55 9.85 13.40 10.55 ;
        RECT  12.90 7.15 13.60 7.85 ;
        RECT  15.80 3.95 16.30 7.85 ;
        RECT  15.60 7.15 16.30 7.85 ;
        RECT  16.85 3.70 17.70 4.45 ;
        RECT  17.20 2.45 17.70 4.45 ;
        RECT  15.80 3.95 17.70 4.45 ;
        RECT  17.20 2.45 17.90 3.15 ;
    END
END NA7X2
MACRO NA7X3
    CLASS CORE ;
    FOREIGN NA7X3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  9.55 7.00 10.75 7.50 ;
        RECT  9.35 2.45 10.05 4.35 ;
        RECT  9.55 2.45 10.05 7.50 ;
        RECT  10.05 7.00 10.75 10.40 ;
        RECT  10.05 8.00 10.95 8.90 ;
        RECT  9.70 9.70 11.45 10.40 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  14.10 5.25 15.15 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.45 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  15.65 9.30 16.55 10.20 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  11.40 8.55 12.80 9.05 ;
        RECT  1.80 7.70 2.50 11.00 ;
        RECT  0.45 10.10 3.85 11.00 ;
        RECT  4.65 7.70 5.35 11.00 ;
        RECT  11.40 7.15 12.10 9.05 ;
        RECT  12.10 8.55 12.80 11.00 ;
        RECT  14.25 7.15 14.95 7.85 ;
        RECT  14.45 7.15 14.95 11.00 ;
        RECT  16.95 7.15 17.75 7.85 ;
        RECT  17.05 7.15 17.75 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.80 2.00 4.50 3.85 ;
        RECT  6.50 2.00 7.20 3.85 ;
        RECT  10.70 2.00 11.40 3.15 ;
        RECT  14.50 2.00 15.20 4.35 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  12.90 7.15 13.75 7.85 ;
        RECT  0.45 6.75 1.15 8.40 ;
        RECT  0.45 2.95 2.25 3.65 ;
        RECT  1.75 2.95 2.25 4.95 ;
        RECT  3.15 6.75 3.85 8.40 ;
        RECT  1.75 4.45 4.90 4.95 ;
        RECT  4.40 4.45 4.90 7.25 ;
        RECT  0.45 6.75 4.90 7.25 ;
        RECT  5.15 3.15 5.85 3.85 ;
        RECT  4.40 5.50 5.80 6.20 ;
        RECT  5.35 3.15 5.85 4.95 ;
        RECT  7.85 3.15 8.55 4.95 ;
        RECT  8.00 3.15 8.50 10.55 ;
        RECT  8.00 3.15 8.55 5.65 ;
        RECT  5.35 4.45 8.55 4.95 ;
        RECT  8.00 7.10 8.70 10.55 ;
        RECT  8.00 4.95 9.10 5.65 ;
        RECT  12.15 3.65 13.40 4.35 ;
        RECT  13.25 3.65 13.40 10.55 ;
        RECT  12.90 3.65 13.40 7.85 ;
        RECT  13.25 7.15 13.75 10.55 ;
        RECT  13.25 9.85 13.95 10.55 ;
        RECT  15.80 3.85 16.30 7.85 ;
        RECT  15.60 7.15 16.30 7.85 ;
        RECT  16.85 3.60 17.70 4.35 ;
        RECT  17.20 2.45 17.70 4.35 ;
        RECT  15.80 3.85 17.70 4.35 ;
        RECT  17.20 2.45 17.90 3.15 ;
    END
END NA7X3
MACRO NA7X4
    CLASS CORE ;
    FOREIGN NA7X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.70 2.75 11.40 4.45 ;
        RECT  10.90 2.75 11.40 6.40 ;
        RECT  10.90 5.90 11.95 6.40 ;
        RECT  11.45 5.90 11.95 10.55 ;
        RECT  11.45 7.15 12.15 10.55 ;
        RECT  11.45 8.00 12.35 8.90 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  15.50 5.25 16.55 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.85 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  17.05 9.30 17.95 10.20 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.40 19.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.70 2.50 11.00 ;
        RECT  0.45 10.10 3.85 11.00 ;
        RECT  4.65 7.70 5.35 11.00 ;
        RECT  10.10 7.15 10.80 11.00 ;
        RECT  12.80 7.15 13.50 11.00 ;
        RECT  15.65 7.15 16.35 11.00 ;
        RECT  18.35 7.15 19.15 7.85 ;
        RECT  18.45 7.15 19.15 11.00 ;
        RECT  0.00 11.00 19.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.80 2.00 4.50 3.85 ;
        RECT  6.50 2.00 7.20 3.85 ;
        RECT  9.35 2.00 10.05 4.45 ;
        RECT  12.05 2.00 12.75 4.45 ;
        RECT  15.90 2.00 16.60 4.45 ;
        RECT  0.00 0.00 19.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 6.75 1.15 8.40 ;
        RECT  0.45 2.95 2.25 3.65 ;
        RECT  1.75 2.95 2.25 4.95 ;
        RECT  3.15 6.75 3.85 8.40 ;
        RECT  1.75 4.45 4.90 4.95 ;
        RECT  4.40 4.45 4.90 7.25 ;
        RECT  0.45 6.75 4.90 7.25 ;
        RECT  5.15 3.15 5.85 3.85 ;
        RECT  4.40 5.50 5.80 6.20 ;
        RECT  5.35 3.15 5.85 4.95 ;
        RECT  7.85 3.15 8.55 4.95 ;
        RECT  8.00 3.15 8.50 10.55 ;
        RECT  8.00 3.15 8.55 5.45 ;
        RECT  5.35 4.45 8.55 4.95 ;
        RECT  8.00 7.10 8.70 10.55 ;
        RECT  8.00 4.95 10.45 5.45 ;
        RECT  9.75 4.95 10.45 5.65 ;
        RECT  13.55 3.75 14.80 4.45 ;
        RECT  14.30 3.75 14.80 10.55 ;
        RECT  13.95 9.85 14.80 10.55 ;
        RECT  14.30 7.15 15.00 7.85 ;
        RECT  17.20 3.95 17.70 7.85 ;
        RECT  17.00 7.15 17.70 7.85 ;
        RECT  18.25 3.70 19.10 4.45 ;
        RECT  18.60 2.45 19.10 4.45 ;
        RECT  17.20 3.95 19.10 4.45 ;
        RECT  18.60 2.45 19.30 3.15 ;
    END
END NA7X4
MACRO NA8X1
    CLASS CORE ;
    FOREIGN NA8X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.75 3.75 11.25 10.55 ;
        RECT  10.75 3.75 11.45 4.45 ;
        RECT  10.75 8.95 12.35 10.55 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  15.50 5.40 16.55 6.30 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  14.25 9.30 15.15 10.20 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  17.05 9.30 17.95 10.20 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.40 19.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.70 2.50 11.00 ;
        RECT  0.45 10.10 3.85 11.00 ;
        RECT  4.65 7.70 5.35 11.00 ;
        RECT  9.50 8.90 10.20 11.00 ;
        RECT  13.05 7.35 13.75 11.00 ;
        RECT  15.75 7.35 16.45 11.00 ;
        RECT  18.45 7.35 19.15 11.00 ;
        RECT  0.00 11.00 19.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.80 2.00 4.50 3.85 ;
        RECT  6.50 2.00 7.20 3.85 ;
        RECT  9.40 2.00 10.10 4.45 ;
        RECT  15.85 2.00 16.55 4.45 ;
        RECT  0.00 0.00 19.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 6.75 1.15 8.40 ;
        RECT  0.45 2.95 2.25 3.65 ;
        RECT  1.75 2.95 2.25 4.95 ;
        RECT  3.15 6.75 3.85 8.40 ;
        RECT  1.75 4.45 4.90 4.95 ;
        RECT  4.40 4.45 4.90 7.25 ;
        RECT  0.45 6.75 4.90 7.25 ;
        RECT  5.15 3.15 5.85 3.85 ;
        RECT  4.40 5.50 5.80 6.20 ;
        RECT  5.35 3.15 5.85 4.95 ;
        RECT  7.85 3.15 8.55 4.95 ;
        RECT  8.00 3.15 8.55 10.55 ;
        RECT  5.35 4.45 8.55 4.95 ;
        RECT  8.00 4.95 8.70 10.55 ;
        RECT  8.00 4.95 10.30 5.65 ;
        RECT  11.10 2.60 12.40 3.30 ;
        RECT  11.90 2.60 12.40 8.05 ;
        RECT  11.70 7.35 12.40 8.05 ;
        RECT  11.90 3.50 13.20 4.20 ;
        RECT  11.90 3.70 14.90 4.20 ;
        RECT  14.40 3.70 14.90 8.05 ;
        RECT  14.40 7.35 15.10 8.05 ;
        RECT  17.30 3.95 17.80 8.05 ;
        RECT  17.10 7.35 17.80 8.05 ;
        RECT  18.20 2.45 18.90 4.45 ;
        RECT  17.30 3.95 18.90 4.45 ;
        RECT  18.20 2.45 19.25 3.15 ;
    END
END NA8X1
MACRO NA8X2
    CLASS CORE ;
    FOREIGN NA8X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.05 6.70 11.20 7.60 ;
        RECT  10.70 2.75 11.20 10.55 ;
        RECT  10.70 2.75 11.40 4.45 ;
        RECT  10.70 8.95 11.55 10.55 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  15.50 5.40 16.55 6.30 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  14.25 9.30 15.15 10.20 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.35 13.75 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  17.05 9.30 17.95 10.20 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.40 19.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.70 2.50 11.00 ;
        RECT  0.45 10.10 3.85 11.00 ;
        RECT  4.65 7.70 5.35 11.00 ;
        RECT  9.50 9.10 10.20 11.00 ;
        RECT  13.05 7.25 13.75 11.00 ;
        RECT  12.20 9.10 13.75 11.00 ;
        RECT  15.75 7.25 16.45 11.00 ;
        RECT  18.45 7.25 19.15 11.00 ;
        RECT  0.00 11.00 19.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.80 2.00 4.50 3.85 ;
        RECT  6.50 2.00 7.20 3.85 ;
        RECT  9.35 2.00 10.05 4.45 ;
        RECT  15.90 2.00 16.60 4.45 ;
        RECT  0.00 0.00 19.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 6.75 1.15 8.40 ;
        RECT  0.45 2.95 2.25 3.65 ;
        RECT  1.75 2.95 2.25 4.95 ;
        RECT  3.15 6.75 3.85 8.40 ;
        RECT  1.75 4.45 4.90 4.95 ;
        RECT  4.40 4.45 4.90 7.25 ;
        RECT  0.45 6.75 4.90 7.25 ;
        RECT  5.15 3.15 5.85 3.85 ;
        RECT  4.40 5.50 5.80 6.20 ;
        RECT  5.35 3.15 5.85 4.95 ;
        RECT  7.85 3.15 8.55 4.95 ;
        RECT  8.00 3.15 8.55 10.55 ;
        RECT  5.35 4.45 8.55 4.95 ;
        RECT  8.00 4.95 8.70 10.55 ;
        RECT  8.00 4.95 10.25 5.65 ;
        RECT  11.85 2.45 12.55 3.15 ;
        RECT  11.90 2.45 12.40 7.95 ;
        RECT  11.70 7.25 12.40 7.95 ;
        RECT  11.90 2.45 12.55 4.50 ;
        RECT  11.90 3.80 13.25 4.50 ;
        RECT  11.90 4.00 14.90 4.50 ;
        RECT  14.40 4.00 14.90 7.95 ;
        RECT  14.40 7.25 15.10 7.95 ;
        RECT  17.30 3.95 17.80 7.95 ;
        RECT  17.10 7.25 17.80 7.95 ;
        RECT  18.25 2.45 18.95 4.45 ;
        RECT  17.30 3.95 18.95 4.45 ;
        RECT  18.25 2.45 19.30 3.15 ;
    END
END NA8X2
MACRO NA8X3
    CLASS CORE ;
    FOREIGN NA8X3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  9.35 2.45 9.40 7.15 ;
        RECT  8.90 4.10 9.40 7.15 ;
        RECT  9.35 2.45 9.85 5.00 ;
        RECT  8.65 4.10 9.85 5.00 ;
        RECT  9.35 2.45 10.05 4.15 ;
        RECT  8.65 4.10 10.05 4.15 ;
        RECT  8.90 6.65 11.25 7.15 ;
        RECT  10.75 6.65 11.25 10.55 ;
        RECT  10.75 8.95 11.55 10.55 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  15.50 5.40 16.55 6.30 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  14.25 9.30 15.15 10.20 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.35 13.75 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  17.05 9.30 17.95 10.20 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.40 19.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.70 2.50 11.00 ;
        RECT  0.45 10.10 3.85 11.00 ;
        RECT  4.65 7.70 5.35 11.00 ;
        RECT  9.50 9.10 10.20 11.00 ;
        RECT  12.20 8.55 12.90 11.00 ;
        RECT  13.05 7.25 13.75 9.05 ;
        RECT  12.20 8.55 13.75 9.05 ;
        RECT  15.75 7.25 16.45 11.00 ;
        RECT  18.45 7.25 19.15 11.00 ;
        RECT  0.00 11.00 19.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.80 2.00 4.50 3.35 ;
        RECT  6.50 2.00 7.20 3.35 ;
        RECT  10.70 2.00 11.40 4.30 ;
        RECT  15.90 2.00 16.60 4.45 ;
        RECT  0.00 0.00 19.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 6.75 1.15 8.40 ;
        RECT  0.45 2.95 2.25 3.65 ;
        RECT  1.75 2.95 2.25 4.95 ;
        RECT  3.15 6.75 3.85 8.40 ;
        RECT  1.75 4.45 4.90 4.95 ;
        RECT  4.40 4.45 4.90 7.25 ;
        RECT  0.45 6.75 4.90 7.25 ;
        RECT  5.15 2.65 5.85 3.35 ;
        RECT  4.40 5.50 5.80 6.20 ;
        RECT  5.35 2.65 5.85 4.30 ;
        RECT  6.85 3.80 7.35 8.10 ;
        RECT  6.85 7.60 8.70 8.10 ;
        RECT  6.85 7.90 9.75 8.10 ;
        RECT  7.70 2.65 8.20 4.30 ;
        RECT  5.35 3.80 8.20 4.30 ;
        RECT  7.70 2.65 8.55 3.35 ;
        RECT  8.00 7.60 8.70 10.55 ;
        RECT  8.00 7.90 9.75 8.60 ;
        RECT  9.85 5.50 10.55 6.20 ;
        RECT  9.85 5.50 12.40 6.00 ;
        RECT  11.90 3.75 12.40 7.95 ;
        RECT  11.70 7.25 12.40 7.95 ;
        RECT  12.55 3.55 13.25 4.25 ;
        RECT  11.90 3.75 14.90 4.25 ;
        RECT  14.40 3.75 14.90 7.95 ;
        RECT  14.40 7.25 15.10 7.95 ;
        RECT  17.30 3.95 17.80 7.95 ;
        RECT  17.10 7.25 17.80 7.95 ;
        RECT  18.25 2.45 18.95 4.45 ;
        RECT  17.30 3.95 18.95 4.45 ;
        RECT  18.25 2.45 19.30 3.15 ;
    END
END NA8X3
MACRO NA8X4
    CLASS CORE ;
    FOREIGN NA8X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.75 2.45 11.55 4.10 ;
        RECT  11.05 2.45 11.55 10.00 ;
        RECT  11.45 2.45 11.55 10.20 ;
        RECT  10.85 7.10 11.55 10.00 ;
        RECT  11.45 9.30 12.35 10.20 ;
        RECT  10.85 9.30 14.35 10.00 ;
        RECT  13.60 9.30 14.35 10.55 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  17.00 5.40 17.95 6.30 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.35 15.15 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  18.45 9.30 19.35 10.20 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.70 2.50 11.00 ;
        RECT  0.45 10.10 3.85 11.00 ;
        RECT  4.65 7.70 5.35 11.00 ;
        RECT  9.50 7.10 10.20 11.00 ;
        RECT  9.50 10.65 12.95 11.00 ;
        RECT  14.45 7.70 15.30 8.40 ;
        RECT  14.80 7.70 15.30 11.00 ;
        RECT  17.15 7.65 17.85 11.00 ;
        RECT  19.85 7.65 20.55 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.80 2.00 4.50 3.35 ;
        RECT  6.50 2.00 7.20 3.35 ;
        RECT  9.40 2.00 10.10 4.10 ;
        RECT  12.10 2.00 12.80 4.10 ;
        RECT  17.30 2.00 18.00 4.45 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 6.75 1.15 8.40 ;
        RECT  0.45 2.95 2.25 3.65 ;
        RECT  1.75 2.95 2.25 4.95 ;
        RECT  3.15 6.75 3.85 8.40 ;
        RECT  1.75 4.45 4.90 4.95 ;
        RECT  4.40 4.45 4.90 7.25 ;
        RECT  0.45 6.75 4.90 7.25 ;
        RECT  5.15 2.65 5.85 3.35 ;
        RECT  4.40 5.50 5.80 6.20 ;
        RECT  5.35 2.65 5.85 4.30 ;
        RECT  5.35 3.80 8.35 4.30 ;
        RECT  8.00 2.65 8.35 10.55 ;
        RECT  7.85 2.65 8.35 5.35 ;
        RECT  8.00 4.85 8.50 10.55 ;
        RECT  7.85 2.65 8.55 3.35 ;
        RECT  8.00 7.15 8.70 10.55 ;
        RECT  7.85 4.85 10.60 5.35 ;
        RECT  9.90 4.85 10.60 5.55 ;
        RECT  13.30 2.45 13.80 8.35 ;
        RECT  13.10 7.65 13.80 8.35 ;
        RECT  13.25 2.45 13.95 3.15 ;
        RECT  13.30 3.80 14.65 4.50 ;
        RECT  13.30 6.75 16.30 7.25 ;
        RECT  15.80 6.75 16.30 8.35 ;
        RECT  15.80 7.65 16.50 8.35 ;
        RECT  18.70 3.95 19.20 8.35 ;
        RECT  18.50 7.65 19.20 8.35 ;
        RECT  19.65 2.45 20.35 4.45 ;
        RECT  18.70 3.95 20.35 4.45 ;
        RECT  19.65 2.45 20.70 3.15 ;
    END
END NA8X4
MACRO NO2I1X1
    CLASS CORE ;
    FOREIGN NO2I1X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.55 7.10 1.25 10.50 ;
        RECT  1.45 2.45 2.15 3.15 ;
        RECT  1.45 2.80 2.55 3.15 ;
        RECT  1.65 2.45 2.15 7.60 ;
        RECT  0.55 7.10 2.15 7.60 ;
        RECT  1.65 2.80 2.55 4.05 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.10 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.90 7.70 3.60 11.00 ;
        RECT  4.45 10.10 5.15 11.00 ;
        RECT  0.00 11.00 5.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.05 2.00 3.75 4.00 ;
        RECT  0.00 0.00 5.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.70 5.50 4.00 6.20 ;
        RECT  3.50 4.45 4.00 7.25 ;
        RECT  3.50 6.75 5.10 7.25 ;
        RECT  4.40 3.30 5.10 4.95 ;
        RECT  3.50 4.45 5.10 4.95 ;
        RECT  4.40 6.75 5.10 8.80 ;
    END
END NO2I1X1
MACRO NO2I1X2
    CLASS CORE ;
    FOREIGN NO2I1X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.15 1.15 10.15 ;
        RECT  1.65 2.80 2.15 7.65 ;
        RECT  0.45 7.15 2.15 7.65 ;
        RECT  1.65 2.80 2.55 4.50 ;
        RECT  0.45 9.45 4.20 10.15 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.48 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 4.10 8.15 5.00 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 7.10 6.55 7.80 ;
        RECT  5.85 7.10 6.55 11.00 ;
        RECT  0.00 11.00 8.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 4.40 ;
        RECT  3.15 2.00 3.85 4.40 ;
        RECT  7.20 2.00 7.90 3.65 ;
        RECT  0.00 0.00 8.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.70 5.50 3.40 6.20 ;
        RECT  5.85 3.00 6.55 3.70 ;
        RECT  6.05 3.00 6.55 6.20 ;
        RECT  2.70 5.70 7.70 6.20 ;
        RECT  7.20 5.70 7.70 8.85 ;
        RECT  7.20 7.10 7.90 8.85 ;
    END
END NO2I1X2
MACRO NO2I1X4
    CLASS CORE ;
    FOREIGN NO2I1X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.15 1.15 9.90 ;
        RECT  1.80 2.45 2.30 7.65 ;
        RECT  0.45 7.15 2.30 7.65 ;
        RECT  1.80 2.45 2.50 5.15 ;
        RECT  4.45 2.50 5.20 5.15 ;
        RECT  1.80 4.65 5.20 5.15 ;
        RECT  4.45 2.80 5.35 3.70 ;
        RECT  0.45 9.20 6.85 9.90 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 7.00 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  10.05 4.10 10.95 5.00 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.95 6.85 9.20 7.55 ;
        RECT  8.50 6.85 9.20 11.00 ;
        RECT  10.00 10.10 10.70 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 4.20 ;
        RECT  3.15 2.00 3.85 4.20 ;
        RECT  5.85 2.00 6.55 4.20 ;
        RECT  10.05 2.00 10.75 3.65 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.60 5.60 4.30 6.30 ;
        RECT  8.70 3.00 9.40 3.70 ;
        RECT  8.90 3.00 9.40 6.30 ;
        RECT  3.60 5.80 10.55 6.30 ;
        RECT  10.05 5.80 10.55 8.85 ;
        RECT  10.05 7.10 10.75 8.85 ;
    END
END NO2I1X4
#MACRO NO2X1
#    CLASS CORE ;
#    FOREIGN NO2X1 0.00 0.00  ;
#    ORIGIN 0.00 0.00 ;
#    SIZE 4.20 BY 13.00 ;
#    SYMMETRY x y r90 ;
#    SITE core ;
#    PIN Q
#        DIRECTION OUTPUT ;
#        ANTENNADIFFAREA 1.0 ;
#        PORT
#        LAYER M1M ;
#        RECT  0.60 7.95 1.30 10.45 ;
#        RECT  1.40 2.90 2.15 3.60 ;
#        RECT  1.65 2.90 2.15 8.90 ;
#        RECT  0.60 7.95 2.15 8.90 ;
#        RECT  1.65 3.80 2.40 4.50 ;
#        RECT  0.60 8.00 2.55 8.90 ;
#        END
#    END Q
#    PIN B
#        DIRECTION INPUT ;
#        ANTENNAGATEAREA 1.75 ;
#        PORT
#        LAYER M1M ;
#        RECT  0.25 4.10 1.15 5.10 ;
#        END
#    END B
#    PIN A
#        DIRECTION INPUT ;
#        ANTENNAGATEAREA 1.75 ;
#        PORT
#        LAYER M1M ;
#        RECT  2.75 5.40 3.95 6.30 ;
#        END
#    END A
#    PIN vdd!
#        DIRECTION INOUT ;
#        USE power ;
#        SHAPE ABUTMENT ;
#        PORT
#        LAYER M1M ;
#        RECT  3.00 7.35 3.70 11.00 ;
#        RECT  0.00 11.00 4.20 13.00 ;
#        END
#    END vdd!
#    PIN gnd!
#        DIRECTION INOUT ;
#        USE ground ;
#        SHAPE ABUTMENT ;
#        PORT
#        LAYER M1M ;
#        RECT  1.40 2.00 2.10 2.25 ;
#        RECT  3.05 2.00 3.75 4.45 ;
#        RECT  0.00 0.00 4.20 2.00 ;
#        END
#    END gnd!
#END NO2X1
MACRO NO2X2
    CLASS CORE ;
    FOREIGN NO2X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.15 1.15 10.15 ;
        RECT  1.65 2.45 2.15 7.65 ;
        RECT  0.45 7.15 2.15 7.65 ;
        RECT  1.65 2.45 2.55 4.05 ;
        RECT  0.45 9.45 4.20 10.15 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.48 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.48 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 7.10 6.55 7.80 ;
        RECT  5.85 7.10 6.55 11.00 ;
        RECT  0.00 11.00 7.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.95 ;
        RECT  3.15 2.00 3.85 3.95 ;
        RECT  4.95 2.00 6.55 3.80 ;
        RECT  0.00 0.00 7.00 2.00 ;
        END
    END gnd!
END NO2X2
MACRO NO2X3
    CLASS CORE ;
    FOREIGN NO2X3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.15 1.15 9.80 ;
        RECT  1.65 2.45 2.15 7.65 ;
        RECT  0.45 7.15 2.15 7.65 ;
        RECT  1.65 2.45 2.55 4.05 ;
        RECT  0.45 9.10 5.55 9.80 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.25 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.25 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.95 6.75 6.45 7.45 ;
        RECT  2.95 6.95 7.95 7.45 ;
        RECT  7.25 6.95 7.95 11.00 ;
        RECT  0.00 11.00 8.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.95 ;
        RECT  3.15 2.00 3.85 3.95 ;
        RECT  4.65 2.00 7.95 3.80 ;
        RECT  0.00 0.00 8.40 2.00 ;
        END
    END gnd!
END NO2X3
MACRO NO2X4
    CLASS CORE ;
    FOREIGN NO2X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.95 2.45 2.45 10.55 ;
        RECT  1.80 2.45 2.55 5.00 ;
        RECT  1.65 4.10 2.55 5.00 ;
        RECT  1.95 7.15 2.65 10.55 ;
        RECT  4.50 2.45 5.20 4.90 ;
        RECT  1.65 4.40 5.20 4.90 ;
        RECT  1.95 9.10 8.40 9.80 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 7.00 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 7.00 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 9.55 1.15 11.00 ;
        RECT  4.45 6.75 9.35 7.45 ;
        RECT  4.45 6.95 10.75 7.45 ;
        RECT  10.05 6.95 10.75 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.95 ;
        RECT  3.15 2.00 3.85 3.95 ;
        RECT  5.85 2.00 6.55 3.95 ;
        RECT  7.35 2.00 10.75 4.70 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
END NO2X4
MACRO NO3I1X1
    CLASS CORE ;
    FOREIGN NO3I1X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.25 6.70 1.15 7.60 ;
        RECT  0.25 7.10 1.65 7.60 ;
        RECT  0.65 4.15 1.15 10.50 ;
        RECT  0.95 2.95 1.15 10.50 ;
        RECT  0.45 6.70 1.15 10.50 ;
        RECT  0.95 2.95 1.65 4.65 ;
        RECT  0.45 7.10 1.65 7.80 ;
        RECT  3.65 2.95 4.35 4.65 ;
        RECT  0.65 4.15 4.35 4.65 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  4.90 7.70 5.60 11.00 ;
        RECT  3.80 10.45 5.60 11.00 ;
        RECT  6.35 10.10 7.95 11.00 ;
        RECT  0.00 11.00 8.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.30 2.00 3.00 3.65 ;
        RECT  5.00 2.00 5.70 3.70 ;
        RECT  0.00 0.00 8.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.90 5.45 2.60 6.15 ;
        RECT  2.10 5.45 2.60 7.25 ;
        RECT  6.35 6.75 7.05 9.10 ;
        RECT  6.35 2.95 7.70 3.65 ;
        RECT  7.20 2.95 7.70 7.25 ;
        RECT  2.10 6.75 7.70 7.25 ;
    END
END NO3I1X1
MACRO NO3I1X2
    CLASS CORE ;
    FOREIGN NO3I1X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.55 7.10 1.25 10.55 ;
        RECT  3.05 5.40 3.95 7.60 ;
        RECT  0.55 7.10 3.95 7.60 ;
        RECT  3.45 2.45 3.95 9.60 ;
        RECT  3.25 5.40 3.95 9.60 ;
        RECT  3.45 2.45 4.15 4.55 ;
        RECT  6.45 2.45 7.15 4.55 ;
        RECT  3.45 4.05 7.15 4.55 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  7.75 5.95 8.45 6.65 ;
        RECT  8.65 5.40 9.55 6.45 ;
        RECT  7.75 5.95 9.55 6.45 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  14.25 4.10 15.15 5.00 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  10.00 8.05 10.70 11.00 ;
        RECT  12.70 7.30 13.40 11.00 ;
        RECT  14.25 10.10 14.95 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.65 2.00 2.25 3.80 ;
        RECT  4.95 2.00 5.65 3.60 ;
        RECT  7.80 2.00 8.50 4.00 ;
        RECT  9.55 2.00 12.05 3.80 ;
        RECT  14.20 2.00 14.90 3.65 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.90 8.05 2.60 10.55 ;
        RECT  4.40 5.00 5.10 5.70 ;
        RECT  4.60 7.10 5.30 10.55 ;
        RECT  1.90 10.05 5.30 10.55 ;
        RECT  5.95 8.05 6.65 10.55 ;
        RECT  4.60 7.10 8.00 7.60 ;
        RECT  7.30 7.10 8.00 9.60 ;
        RECT  7.70 4.45 8.20 5.50 ;
        RECT  4.40 5.00 8.20 5.50 ;
        RECT  8.65 7.10 9.35 10.55 ;
        RECT  5.95 10.05 9.35 10.55 ;
        RECT  8.65 7.10 12.05 7.60 ;
        RECT  11.35 7.10 12.05 10.55 ;
        RECT  12.85 2.95 13.55 3.65 ;
        RECT  7.70 4.45 13.55 4.95 ;
        RECT  13.05 2.95 13.55 6.05 ;
        RECT  13.05 5.55 14.70 6.05 ;
        RECT  14.20 5.55 14.70 8.85 ;
        RECT  14.20 7.15 14.90 8.85 ;
    END
END NO3I1X2
MACRO NO3I1X4
    CLASS CORE ;
    FOREIGN NO3I1X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.85 6.35 6.95 6.70 ;
        RECT  0.85 6.20 1.55 10.55 ;
        RECT  3.55 6.20 4.25 9.60 ;
        RECT  5.85 5.40 6.75 6.70 ;
        RECT  6.25 2.50 6.75 9.60 ;
        RECT  0.85 6.20 6.75 6.70 ;
        RECT  6.25 2.50 6.95 4.75 ;
        RECT  6.25 6.35 6.95 9.60 ;
        RECT  8.95 2.50 9.65 4.75 ;
        RECT  11.65 2.50 12.35 4.75 ;
        RECT  6.25 4.25 12.35 4.75 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.30 16.55 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  13.90 5.30 15.15 6.30 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  22.65 4.10 23.55 5.00 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  15.70 7.70 16.40 11.00 ;
        RECT  18.40 7.70 19.10 11.00 ;
        RECT  21.10 7.30 21.80 11.00 ;
        RECT  22.65 10.10 23.35 11.00 ;
        RECT  0.00 11.00 23.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.70 2.00 4.10 3.80 ;
        RECT  4.90 2.00 5.60 3.65 ;
        RECT  7.60 2.00 8.30 3.65 ;
        RECT  10.30 2.00 11.00 3.65 ;
        RECT  13.00 2.00 13.70 3.65 ;
        RECT  15.15 2.00 20.35 3.80 ;
        RECT  22.60 2.00 23.30 3.65 ;
        RECT  0.00 0.00 23.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.20 7.15 2.90 10.55 ;
        RECT  4.90 7.15 5.60 10.55 ;
        RECT  7.20 5.20 7.90 5.90 ;
        RECT  7.60 6.75 8.30 10.55 ;
        RECT  2.20 10.05 8.30 10.55 ;
        RECT  8.95 7.70 9.65 10.55 ;
        RECT  10.30 6.75 11.00 9.60 ;
        RECT  11.65 7.70 12.35 10.55 ;
        RECT  7.60 6.75 13.70 7.25 ;
        RECT  12.95 4.35 13.45 5.70 ;
        RECT  7.20 5.20 13.45 5.70 ;
        RECT  13.00 6.75 13.70 9.60 ;
        RECT  14.35 6.75 15.05 10.55 ;
        RECT  8.95 10.05 15.05 10.55 ;
        RECT  17.05 6.75 17.75 10.55 ;
        RECT  14.35 6.75 20.45 7.25 ;
        RECT  19.75 6.75 20.45 10.55 ;
        RECT  21.25 2.95 21.95 3.65 ;
        RECT  12.95 4.35 21.95 4.85 ;
        RECT  21.45 2.95 21.95 6.05 ;
        RECT  21.45 5.55 23.10 6.05 ;
        RECT  22.60 5.55 23.10 8.90 ;
        RECT  22.60 7.30 23.30 8.90 ;
    END
END NO3I1X4
MACRO NO3I2X1
    CLASS CORE ;
    FOREIGN NO3I2X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.65 4.45 7.60 ;
        RECT  3.75 2.45 3.90 10.50 ;
        RECT  3.20 2.45 3.90 4.05 ;
        RECT  3.75 3.55 4.25 10.50 ;
        RECT  3.75 6.65 4.45 10.50 ;
        RECT  5.90 2.45 6.60 4.05 ;
        RECT  3.20 3.55 6.60 4.05 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.30 6.75 6.30 ;
        RECT  5.85 5.30 7.25 6.00 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.40 9.55 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.55 7.20 1.25 11.00 ;
        RECT  0.45 10.10 2.95 11.00 ;
        RECT  7.10 7.70 7.80 11.00 ;
        RECT  8.65 10.10 9.35 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.65 2.00 2.35 2.40 ;
        RECT  4.55 2.00 5.25 3.10 ;
        RECT  7.25 2.00 7.95 3.10 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.65 3.05 2.40 3.75 ;
        RECT  1.90 3.05 2.40 8.80 ;
        RECT  1.90 7.20 2.60 8.80 ;
        RECT  1.90 5.30 3.30 6.00 ;
        RECT  4.70 4.50 5.40 5.20 ;
        RECT  4.90 4.50 5.40 7.25 ;
        RECT  7.70 3.55 8.20 7.25 ;
        RECT  4.90 6.75 9.10 7.25 ;
        RECT  8.60 2.45 9.10 4.05 ;
        RECT  7.70 3.55 9.10 4.05 ;
        RECT  8.60 6.75 9.10 9.10 ;
        RECT  8.60 2.45 9.30 3.15 ;
        RECT  8.60 7.50 9.30 9.10 ;
    END
END NO3I2X1
MACRO NO3I2X2
    CLASS CORE ;
    FOREIGN NO3I2X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  3.35 7.10 4.05 10.55 ;
        RECT  5.85 5.40 6.75 7.60 ;
        RECT  3.35 7.10 6.75 7.60 ;
        RECT  6.25 2.45 6.75 9.60 ;
        RECT  6.05 5.40 6.75 9.60 ;
        RECT  6.25 2.45 6.95 4.55 ;
        RECT  9.25 2.45 9.95 4.55 ;
        RECT  6.25 4.05 9.95 4.55 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  17.05 4.10 17.95 5.00 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 7.15 1.20 11.00 ;
        RECT  0.50 10.10 2.40 11.00 ;
        RECT  12.80 8.05 13.50 11.00 ;
        RECT  15.50 7.30 16.20 11.00 ;
        RECT  17.05 10.10 17.75 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 2.00 1.20 4.05 ;
        RECT  3.35 2.00 4.95 3.80 ;
        RECT  7.75 2.00 8.45 3.60 ;
        RECT  10.60 2.00 11.30 4.00 ;
        RECT  12.35 2.00 14.85 3.80 ;
        RECT  17.00 2.00 17.70 3.65 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.85 3.35 2.55 4.05 ;
        RECT  2.05 3.35 2.55 8.85 ;
        RECT  1.85 7.15 2.55 8.85 ;
        RECT  2.05 5.95 4.95 6.45 ;
        RECT  4.25 5.95 4.95 6.65 ;
        RECT  4.70 8.05 5.40 10.55 ;
        RECT  7.40 7.10 8.10 10.55 ;
        RECT  4.70 10.05 8.10 10.55 ;
        RECT  8.75 8.05 9.45 10.55 ;
        RECT  7.40 7.10 10.80 7.60 ;
        RECT  10.10 7.10 10.80 9.60 ;
        RECT  10.75 4.45 11.25 6.65 ;
        RECT  10.55 5.95 11.25 6.65 ;
        RECT  11.45 7.10 12.15 10.55 ;
        RECT  8.75 10.05 12.15 10.55 ;
        RECT  11.45 7.10 14.85 7.60 ;
        RECT  14.15 7.10 14.85 10.55 ;
        RECT  15.65 2.95 16.35 3.65 ;
        RECT  10.75 4.45 16.35 4.95 ;
        RECT  15.85 2.95 16.35 6.05 ;
        RECT  15.85 5.55 17.50 6.05 ;
        RECT  17.00 5.55 17.50 8.85 ;
        RECT  17.00 7.15 17.70 8.85 ;
    END
END NO3I2X2
MACRO NO3I2X4
    CLASS CORE ;
    FOREIGN NO3I2X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 26.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  3.65 6.20 4.35 10.55 ;
        RECT  6.35 6.20 7.05 9.60 ;
        RECT  3.65 6.20 9.75 6.70 ;
        RECT  9.05 2.50 9.55 9.60 ;
        RECT  8.65 5.40 9.55 6.70 ;
        RECT  9.05 2.50 9.75 4.75 ;
        RECT  9.05 6.20 9.75 9.60 ;
        RECT  11.75 2.50 12.45 4.75 ;
        RECT  14.45 2.50 15.15 4.75 ;
        RECT  9.05 4.25 15.15 4.75 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.30 19.35 6.30 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  25.45 4.10 26.35 5.00 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.20 1.15 11.00 ;
        RECT  0.45 10.10 2.40 11.00 ;
        RECT  18.50 7.70 19.20 11.00 ;
        RECT  21.20 7.70 21.90 11.00 ;
        RECT  23.90 7.30 24.60 11.00 ;
        RECT  25.45 10.10 26.15 11.00 ;
        RECT  0.00 11.00 26.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.65 ;
        RECT  3.30 2.00 6.85 3.80 ;
        RECT  7.70 2.00 8.40 3.65 ;
        RECT  10.40 2.00 11.10 3.65 ;
        RECT  13.10 2.00 13.80 3.65 ;
        RECT  15.80 2.00 16.50 3.65 ;
        RECT  17.35 2.00 22.55 3.80 ;
        RECT  25.40 2.00 26.10 3.65 ;
        RECT  0.00 0.00 26.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 2.95 2.30 8.80 ;
        RECT  1.80 2.95 2.50 3.65 ;
        RECT  1.80 7.20 2.50 8.80 ;
        RECT  5.00 7.15 5.70 10.55 ;
        RECT  1.80 5.05 8.10 5.55 ;
        RECT  7.40 5.05 8.10 5.75 ;
        RECT  7.70 7.15 8.40 10.55 ;
        RECT  10.40 6.75 11.10 10.55 ;
        RECT  5.00 10.05 11.10 10.55 ;
        RECT  11.75 7.70 12.45 10.55 ;
        RECT  12.65 5.20 13.35 5.90 ;
        RECT  13.10 6.75 13.80 9.60 ;
        RECT  14.45 7.70 15.15 10.55 ;
        RECT  10.40 6.75 16.50 7.25 ;
        RECT  15.80 6.75 16.50 9.60 ;
        RECT  16.45 4.35 16.95 5.70 ;
        RECT  12.65 5.20 16.95 5.70 ;
        RECT  17.15 6.75 17.85 10.55 ;
        RECT  11.75 10.05 17.85 10.55 ;
        RECT  19.85 6.75 20.55 10.55 ;
        RECT  17.15 6.75 23.25 7.25 ;
        RECT  22.55 6.75 23.25 10.55 ;
        RECT  24.05 2.95 24.75 3.65 ;
        RECT  16.45 4.35 24.75 4.85 ;
        RECT  24.25 2.95 24.75 6.05 ;
        RECT  24.25 5.55 25.90 6.05 ;
        RECT  25.40 5.55 25.90 8.90 ;
        RECT  25.40 7.30 26.10 8.90 ;
    END
END NO3I2X4
MACRO NO3X1
    CLASS CORE ;
    FOREIGN NO3X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.10 1.15 9.75 ;
        RECT  1.65 6.65 2.95 7.80 ;
        RECT  2.45 4.15 2.95 7.80 ;
        RECT  0.45 7.10 2.95 7.80 ;
        RECT  3.15 2.95 3.85 4.65 ;
        RECT  5.85 3.00 6.55 4.65 ;
        RECT  2.45 4.15 6.55 4.65 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.90 5.25 5.35 5.95 ;
        RECT  4.45 5.25 5.35 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.35 1.15 6.35 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  5.80 7.70 6.50 11.00 ;
        RECT  0.00 11.00 7.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 3.65 ;
        RECT  4.50 2.00 5.20 3.65 ;
        RECT  0.00 0.00 7.00 2.00 ;
        END
    END gnd!
END NO3X1
MACRO NO3X2
    CLASS CORE ;
    FOREIGN NO3X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.55 6.75 1.25 10.55 ;
        RECT  2.05 4.45 2.55 7.25 ;
        RECT  1.65 5.40 2.55 7.25 ;
        RECT  0.55 6.75 3.95 7.25 ;
        RECT  3.25 6.75 3.95 9.60 ;
        RECT  5.45 2.45 6.15 4.95 ;
        RECT  8.15 2.45 8.85 4.95 ;
        RECT  2.05 4.45 8.85 4.95 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  10.00 7.70 10.70 11.00 ;
        RECT  12.70 7.30 13.40 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 3.05 3.80 ;
        RECT  4.10 2.00 4.80 4.00 ;
        RECT  6.80 2.00 7.50 4.00 ;
        RECT  9.95 2.00 13.55 3.80 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.90 7.70 2.60 10.55 ;
        RECT  4.60 6.75 5.30 10.55 ;
        RECT  1.90 10.05 5.30 10.55 ;
        RECT  5.95 7.70 6.65 10.55 ;
        RECT  4.60 6.75 8.00 7.25 ;
        RECT  7.30 6.75 8.00 9.60 ;
        RECT  8.65 6.75 9.35 10.55 ;
        RECT  5.95 10.05 9.35 10.55 ;
        RECT  8.65 6.75 12.05 7.25 ;
        RECT  11.35 6.75 12.05 10.55 ;
    END
END NO3X2
MACRO NO3X3
    CLASS CORE ;
    FOREIGN NO3X3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.95 5.85 2.65 10.55 ;
        RECT  3.50 3.15 4.00 6.35 ;
        RECT  3.05 5.40 4.00 6.35 ;
        RECT  1.95 5.85 5.35 6.35 ;
        RECT  4.65 5.85 5.35 9.60 ;
        RECT  5.30 2.45 6.00 3.65 ;
        RECT  8.00 2.45 8.70 3.65 ;
        RECT  10.70 2.45 11.40 3.65 ;
        RECT  3.50 3.15 11.40 3.65 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 7.35 ;
        PORT
        LAYER M1M ;
        RECT  11.45 4.10 12.35 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 7.35 ;
        PORT
        LAYER M1M ;
        RECT  7.25 4.10 8.15 5.00 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 7.35 ;
        PORT
        LAYER M1M ;
        RECT  4.45 4.10 5.35 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 9.55 1.15 11.00 ;
        RECT  11.40 6.80 12.10 11.00 ;
        RECT  14.10 6.80 14.80 11.00 ;
        RECT  15.65 9.55 16.35 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 3.05 3.80 ;
        RECT  3.95 2.00 4.65 2.70 ;
        RECT  6.65 2.00 7.35 2.70 ;
        RECT  9.35 2.00 10.05 2.70 ;
        RECT  12.05 2.00 12.75 2.70 ;
        RECT  13.65 2.00 16.35 3.80 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.30 6.80 4.00 10.55 ;
        RECT  6.00 5.85 6.70 10.55 ;
        RECT  3.30 10.05 6.70 10.55 ;
        RECT  7.35 6.80 8.05 10.55 ;
        RECT  6.00 5.85 9.40 6.35 ;
        RECT  8.70 5.85 9.40 9.60 ;
        RECT  10.05 5.85 10.75 10.55 ;
        RECT  7.35 10.05 10.75 10.55 ;
        RECT  10.05 5.85 13.45 6.35 ;
        RECT  12.75 5.85 13.45 10.55 ;
    END
END NO3X3
MACRO NO3X4
    CLASS CORE ;
    FOREIGN NO3X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  3.30 5.85 4.00 9.60 ;
        RECT  5.85 5.40 6.70 6.35 ;
        RECT  3.30 5.85 6.70 6.35 ;
        RECT  6.30 3.15 6.70 9.60 ;
        RECT  6.00 5.40 6.70 9.60 ;
        RECT  6.30 3.15 6.80 6.30 ;
        RECT  3.30 5.85 6.80 6.30 ;
        RECT  9.60 2.45 10.30 3.65 ;
        RECT  12.30 2.45 13.00 3.65 ;
        RECT  15.00 2.45 15.70 3.65 ;
        RECT  6.30 3.15 15.70 3.65 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  15.65 4.10 16.55 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  11.45 4.10 12.35 5.00 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.55 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 9.55 1.15 11.00 ;
        RECT  15.75 6.80 16.45 11.00 ;
        RECT  18.45 6.80 19.15 11.00 ;
        RECT  21.15 6.80 21.85 11.00 ;
        RECT  22.65 9.55 23.35 11.00 ;
        RECT  0.00 11.00 23.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 5.65 3.80 ;
        RECT  8.25 2.00 8.95 2.70 ;
        RECT  10.95 2.00 11.65 2.70 ;
        RECT  13.65 2.00 14.35 2.70 ;
        RECT  16.35 2.00 17.05 2.70 ;
        RECT  17.95 2.00 23.35 3.80 ;
        RECT  0.00 0.00 23.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.95 6.80 2.65 10.55 ;
        RECT  4.65 6.80 5.35 10.55 ;
        RECT  7.35 5.85 8.05 10.55 ;
        RECT  1.95 10.05 8.05 10.55 ;
        RECT  8.85 6.80 9.55 10.55 ;
        RECT  10.20 5.85 10.90 9.60 ;
        RECT  11.55 6.80 12.25 10.55 ;
        RECT  7.35 5.85 13.60 6.35 ;
        RECT  12.90 5.85 13.60 9.60 ;
        RECT  14.25 5.85 14.95 10.55 ;
        RECT  8.85 10.05 14.95 10.55 ;
        RECT  17.10 5.85 17.80 10.55 ;
        RECT  14.25 5.85 20.50 6.35 ;
        RECT  19.80 5.85 20.50 10.55 ;
    END
END NO3X4
MACRO NO4I1X1
    CLASS CORE ;
    FOREIGN NO4I1X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  14.25 2.80 14.75 8.75 ;
        RECT  14.05 7.10 14.75 8.75 ;
        RECT  14.25 2.80 15.15 3.70 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  12.35 5.40 13.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  10.05 4.10 10.95 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 3.95 5.00 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.15 1.15 11.00 ;
        RECT  0.45 10.10 2.50 11.00 ;
        RECT  5.80 8.55 6.50 11.00 ;
        RECT  8.80 7.55 9.50 11.00 ;
        RECT  12.70 7.30 13.40 11.00 ;
        RECT  12.70 10.10 14.95 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.75 2.00 3.45 3.20 ;
        RECT  5.45 2.00 6.15 3.20 ;
        RECT  5.65 2.00 6.15 4.80 ;
        RECT  5.65 4.10 6.85 4.80 ;
        RECT  7.75 2.00 9.35 2.90 ;
        RECT  10.20 2.00 10.90 3.65 ;
        RECT  12.90 2.00 13.60 3.70 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  7.30 7.55 8.00 8.25 ;
        RECT  1.40 2.55 2.30 3.25 ;
        RECT  1.80 2.55 2.30 8.85 ;
        RECT  1.80 6.65 2.50 8.85 ;
        RECT  3.30 7.60 4.00 10.10 ;
        RECT  4.10 2.55 4.90 3.25 ;
        RECT  4.40 2.55 4.90 5.85 ;
        RECT  5.00 6.45 5.70 7.15 ;
        RECT  1.80 6.65 5.70 7.15 ;
        RECT  4.40 5.35 6.85 5.85 ;
        RECT  6.15 5.35 6.65 8.10 ;
        RECT  3.30 7.60 6.65 8.10 ;
        RECT  6.15 5.35 6.85 6.05 ;
        RECT  7.50 4.35 7.80 10.55 ;
        RECT  7.30 4.35 7.80 8.25 ;
        RECT  7.50 7.55 8.00 10.55 ;
        RECT  7.50 9.85 8.20 10.55 ;
        RECT  8.25 5.35 8.95 6.05 ;
        RECT  8.50 4.10 9.20 4.85 ;
        RECT  7.30 4.35 9.20 4.85 ;
        RECT  11.40 2.95 11.70 10.05 ;
        RECT  11.15 5.55 11.70 10.05 ;
        RECT  11.15 7.55 11.85 10.05 ;
        RECT  11.40 2.95 11.90 6.05 ;
        RECT  8.25 5.55 11.90 6.05 ;
        RECT  11.40 2.95 12.25 3.65 ;
    END
END NO4I1X1
MACRO NO4I1X2
    CLASS CORE ;
    FOREIGN NO4I1X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  14.25 2.45 14.75 10.50 ;
        RECT  14.05 7.10 14.75 10.50 ;
        RECT  14.25 2.45 15.15 4.10 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  12.35 5.40 13.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  10.05 4.10 10.95 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 3.95 5.00 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.15 1.15 11.00 ;
        RECT  0.45 10.10 2.50 11.00 ;
        RECT  5.80 8.55 6.50 11.00 ;
        RECT  8.80 7.55 9.50 11.00 ;
        RECT  12.70 7.30 13.40 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.75 2.00 3.45 3.20 ;
        RECT  5.45 2.00 6.15 3.20 ;
        RECT  5.65 2.00 6.15 4.80 ;
        RECT  5.65 4.10 6.85 4.80 ;
        RECT  7.65 2.00 9.25 2.90 ;
        RECT  10.05 2.00 10.75 3.15 ;
        RECT  12.90 2.00 13.60 4.10 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  7.30 7.55 8.00 8.25 ;
        RECT  1.40 2.55 2.30 3.25 ;
        RECT  1.80 2.55 2.30 8.85 ;
        RECT  1.80 6.65 2.50 8.85 ;
        RECT  3.30 7.60 4.00 10.10 ;
        RECT  4.10 2.55 4.90 3.25 ;
        RECT  4.40 2.55 4.90 5.85 ;
        RECT  5.00 6.45 5.70 7.15 ;
        RECT  1.80 6.65 5.70 7.15 ;
        RECT  4.40 5.35 6.85 5.85 ;
        RECT  6.15 5.35 6.65 8.10 ;
        RECT  3.30 7.60 6.65 8.10 ;
        RECT  6.15 5.35 6.85 6.05 ;
        RECT  7.50 4.35 7.80 10.55 ;
        RECT  7.30 4.35 7.80 8.25 ;
        RECT  7.50 7.55 8.00 10.55 ;
        RECT  7.50 9.85 8.20 10.55 ;
        RECT  8.25 5.35 8.95 6.05 ;
        RECT  8.50 4.10 9.20 4.85 ;
        RECT  7.30 4.35 9.20 4.85 ;
        RECT  11.40 2.45 11.70 10.05 ;
        RECT  11.15 5.55 11.70 10.05 ;
        RECT  11.15 7.55 11.85 10.05 ;
        RECT  11.40 2.45 11.90 6.05 ;
        RECT  8.25 5.55 11.90 6.05 ;
        RECT  11.40 2.45 12.10 3.15 ;
    END
END NO4I1X2
MACRO NO4I1X4
    CLASS CORE ;
    FOREIGN NO4I1X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  14.25 2.45 14.75 10.50 ;
        RECT  14.05 7.10 14.75 10.50 ;
        RECT  14.25 2.45 14.95 4.10 ;
        RECT  14.25 5.35 15.15 6.30 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  12.35 5.40 13.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  10.05 4.10 10.95 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 3.95 5.00 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.15 1.15 11.00 ;
        RECT  0.45 10.10 2.50 11.00 ;
        RECT  5.80 8.55 6.50 11.00 ;
        RECT  8.80 7.55 9.50 11.00 ;
        RECT  12.70 7.30 13.40 11.00 ;
        RECT  15.40 7.30 16.10 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.75 2.00 3.45 3.20 ;
        RECT  5.45 2.00 6.15 3.20 ;
        RECT  5.65 2.00 6.15 4.80 ;
        RECT  5.65 4.10 6.85 4.80 ;
        RECT  7.15 2.00 8.75 2.90 ;
        RECT  10.05 2.00 10.75 3.15 ;
        RECT  12.90 2.00 13.60 4.10 ;
        RECT  15.60 2.00 16.30 4.10 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  7.30 7.55 8.00 8.25 ;
        RECT  1.40 2.55 2.30 3.25 ;
        RECT  1.80 2.55 2.30 8.85 ;
        RECT  1.80 6.65 2.50 8.85 ;
        RECT  3.30 7.60 4.00 10.10 ;
        RECT  4.10 2.55 4.90 3.25 ;
        RECT  4.40 2.55 4.90 5.85 ;
        RECT  5.00 6.45 5.70 7.15 ;
        RECT  1.80 6.65 5.70 7.15 ;
        RECT  4.40 5.35 6.85 5.85 ;
        RECT  6.15 5.35 6.65 8.10 ;
        RECT  3.30 7.60 6.65 8.10 ;
        RECT  6.15 5.35 6.85 6.05 ;
        RECT  7.50 4.35 7.80 10.55 ;
        RECT  7.30 4.35 7.80 8.25 ;
        RECT  7.50 7.55 8.00 10.55 ;
        RECT  7.50 9.85 8.20 10.55 ;
        RECT  8.25 5.35 8.95 6.05 ;
        RECT  8.50 4.10 9.20 4.85 ;
        RECT  7.30 4.35 9.20 4.85 ;
        RECT  11.40 2.45 11.70 10.05 ;
        RECT  11.15 5.55 11.70 10.05 ;
        RECT  11.15 7.55 11.85 10.05 ;
        RECT  11.40 2.45 11.90 6.05 ;
        RECT  8.25 5.55 11.90 6.05 ;
        RECT  11.40 2.45 12.10 3.15 ;
    END
END NO4I1X4
MACRO NO4I2X1
    CLASS CORE ;
    FOREIGN NO4I2X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  12.85 2.80 13.35 8.70 ;
        RECT  12.85 7.10 13.55 8.70 ;
        RECT  12.85 2.80 13.75 3.70 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  10.95 5.40 12.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.55 5.00 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 3.05 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.90 2.50 11.00 ;
        RECT  4.65 7.90 5.35 11.00 ;
        RECT  3.45 10.10 6.05 11.00 ;
        RECT  7.65 7.55 8.35 11.00 ;
        RECT  11.50 7.30 12.20 11.00 ;
        RECT  11.50 10.10 13.55 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.15 2.00 2.85 4.25 ;
        RECT  2.00 3.55 2.85 4.25 ;
        RECT  4.80 4.10 5.50 4.80 ;
        RECT  6.15 2.00 6.65 4.60 ;
        RECT  4.80 4.10 6.65 4.60 ;
        RECT  6.15 2.00 7.95 2.90 ;
        RECT  8.80 2.00 9.50 3.60 ;
        RECT  11.50 2.00 12.20 3.65 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.30 2.45 0.80 9.55 ;
        RECT  0.30 2.45 1.00 4.25 ;
        RECT  0.30 7.95 1.15 9.55 ;
        RECT  0.30 3.55 1.35 4.25 ;
        RECT  1.25 6.75 1.95 7.45 ;
        RECT  1.25 6.75 4.00 7.25 ;
        RECT  3.50 2.50 4.00 8.55 ;
        RECT  3.30 6.75 4.00 8.55 ;
        RECT  3.50 2.50 5.20 3.20 ;
        RECT  6.15 7.85 7.00 8.55 ;
        RECT  6.50 5.45 6.85 10.55 ;
        RECT  6.35 5.45 6.85 8.55 ;
        RECT  6.50 7.85 7.00 10.55 ;
        RECT  6.50 9.85 7.20 10.55 ;
        RECT  7.15 4.10 7.65 5.95 ;
        RECT  6.35 5.45 7.65 5.95 ;
        RECT  7.15 4.10 7.85 4.85 ;
        RECT  7.30 6.40 8.00 7.10 ;
        RECT  7.30 6.60 10.50 7.10 ;
        RECT  10.00 2.90 10.50 10.45 ;
        RECT  10.00 7.55 10.70 10.45 ;
        RECT  10.00 2.90 10.85 3.60 ;
    END
END NO4I2X1
MACRO NO4I2X2
    CLASS CORE ;
    FOREIGN NO4I2X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  12.85 2.45 13.35 10.50 ;
        RECT  12.85 7.10 13.55 10.50 ;
        RECT  12.85 2.45 13.75 4.10 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  10.95 5.40 12.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.55 5.00 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 3.05 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.90 2.50 11.00 ;
        RECT  4.65 7.90 5.35 11.00 ;
        RECT  3.45 10.10 6.05 11.00 ;
        RECT  7.65 7.55 8.35 11.00 ;
        RECT  11.50 7.30 12.20 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.15 2.00 2.85 4.25 ;
        RECT  2.00 3.55 2.85 4.25 ;
        RECT  4.80 4.10 5.50 4.80 ;
        RECT  6.15 2.00 6.65 4.60 ;
        RECT  4.80 4.10 6.65 4.60 ;
        RECT  6.15 2.00 7.05 2.90 ;
        RECT  8.65 2.00 9.35 3.15 ;
        RECT  11.50 2.00 12.20 4.10 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.30 2.45 0.80 9.55 ;
        RECT  0.30 2.45 1.00 4.25 ;
        RECT  0.30 7.95 1.15 9.55 ;
        RECT  0.30 3.55 1.35 4.25 ;
        RECT  1.25 6.75 1.95 7.45 ;
        RECT  1.25 6.75 4.00 7.25 ;
        RECT  3.50 2.50 4.00 8.50 ;
        RECT  3.30 6.75 4.00 8.50 ;
        RECT  3.50 2.50 5.20 3.20 ;
        RECT  6.15 7.85 7.00 8.55 ;
        RECT  6.50 5.45 6.75 10.55 ;
        RECT  6.25 5.45 6.75 8.55 ;
        RECT  6.50 7.85 7.00 10.55 ;
        RECT  6.50 9.85 7.20 10.55 ;
        RECT  7.15 4.10 7.65 5.95 ;
        RECT  6.25 5.45 7.65 5.95 ;
        RECT  7.15 4.10 7.85 4.85 ;
        RECT  7.20 6.40 7.90 7.10 ;
        RECT  7.20 6.60 10.50 7.10 ;
        RECT  10.00 2.45 10.50 10.45 ;
        RECT  10.00 2.45 10.70 3.15 ;
        RECT  10.00 7.55 10.70 10.45 ;
    END
END NO4I2X2
MACRO NO4I2X4
    CLASS CORE ;
    FOREIGN NO4I2X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  12.85 2.75 13.35 10.50 ;
        RECT  12.85 2.75 13.55 4.35 ;
        RECT  12.85 7.10 13.55 10.50 ;
        RECT  12.85 8.00 13.75 8.90 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  10.95 5.40 12.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.55 5.00 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 3.05 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.90 2.50 11.00 ;
        RECT  4.65 7.90 5.35 11.00 ;
        RECT  3.45 10.10 6.05 11.00 ;
        RECT  7.65 7.55 8.35 11.00 ;
        RECT  11.50 7.30 12.20 11.00 ;
        RECT  14.20 7.30 14.90 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.15 2.00 2.85 4.25 ;
        RECT  2.00 3.55 2.85 4.25 ;
        RECT  4.80 4.10 5.50 4.80 ;
        RECT  6.15 2.00 6.65 4.60 ;
        RECT  4.80 4.10 6.65 4.60 ;
        RECT  6.15 2.00 7.20 2.90 ;
        RECT  8.65 2.00 9.35 3.45 ;
        RECT  11.50 2.00 12.20 4.40 ;
        RECT  14.20 2.00 14.90 4.40 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.30 2.45 0.80 9.55 ;
        RECT  0.30 2.45 1.00 4.25 ;
        RECT  0.30 7.95 1.15 9.55 ;
        RECT  0.30 3.55 1.35 4.25 ;
        RECT  1.25 6.75 1.95 7.45 ;
        RECT  1.25 6.75 4.00 7.25 ;
        RECT  3.50 2.50 4.00 8.50 ;
        RECT  3.30 6.75 4.00 8.50 ;
        RECT  3.50 2.50 5.20 3.20 ;
        RECT  6.15 7.85 7.00 8.55 ;
        RECT  6.50 5.45 6.75 10.55 ;
        RECT  6.25 5.45 6.75 8.55 ;
        RECT  6.50 7.85 7.00 10.55 ;
        RECT  6.50 9.85 7.20 10.55 ;
        RECT  7.15 4.10 7.65 5.95 ;
        RECT  6.25 5.45 7.65 5.95 ;
        RECT  7.15 4.10 7.85 4.85 ;
        RECT  7.20 6.40 7.90 7.10 ;
        RECT  7.20 6.60 10.50 7.10 ;
        RECT  10.00 2.75 10.50 10.45 ;
        RECT  10.00 2.75 10.70 3.45 ;
        RECT  10.00 7.55 10.70 10.45 ;
    END
END NO4I2X4
MACRO NO4I3X1
    CLASS CORE ;
    FOREIGN NO4I3X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  14.25 2.80 14.75 8.70 ;
        RECT  14.25 7.10 14.95 8.70 ;
        RECT  14.25 2.80 15.15 4.20 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  9.55 5.40 10.95 6.15 ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  12.50 5.40 13.75 6.30 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 3.05 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.90 2.50 11.00 ;
        RECT  4.65 7.90 5.35 11.00 ;
        RECT  3.30 10.10 5.90 11.00 ;
        RECT  7.50 7.70 8.20 11.00 ;
        RECT  12.90 7.30 13.60 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.15 2.00 2.85 4.25 ;
        RECT  2.00 3.55 2.85 4.25 ;
        RECT  4.80 4.10 5.50 4.80 ;
        RECT  6.05 2.00 6.55 4.60 ;
        RECT  4.80 4.10 6.55 4.60 ;
        RECT  7.15 2.00 7.85 3.10 ;
        RECT  9.85 2.00 10.55 3.10 ;
        RECT  12.90 2.00 13.60 4.20 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.30 2.45 0.80 9.55 ;
        RECT  0.30 2.45 1.00 4.25 ;
        RECT  0.30 7.95 1.15 9.55 ;
        RECT  0.30 3.55 1.35 4.25 ;
        RECT  1.25 6.75 1.95 7.45 ;
        RECT  1.25 6.75 4.00 7.25 ;
        RECT  3.50 2.50 4.00 8.50 ;
        RECT  3.30 6.75 4.00 8.50 ;
        RECT  3.50 2.50 5.20 3.20 ;
        RECT  6.00 7.85 6.85 8.55 ;
        RECT  6.35 5.45 6.70 10.55 ;
        RECT  6.20 5.45 6.70 8.55 ;
        RECT  6.35 7.85 6.85 10.55 ;
        RECT  6.35 9.85 7.05 10.55 ;
        RECT  7.15 4.10 7.65 5.95 ;
        RECT  6.20 5.45 7.65 5.95 ;
        RECT  7.15 4.10 7.85 4.85 ;
        RECT  7.15 6.40 7.85 7.25 ;
        RECT  8.50 2.45 9.00 7.25 ;
        RECT  8.50 2.45 9.20 3.15 ;
        RECT  7.15 6.75 10.35 7.25 ;
        RECT  9.85 6.75 10.35 10.45 ;
        RECT  9.85 7.55 10.55 10.45 ;
        RECT  11.05 2.45 12.05 3.15 ;
        RECT  11.55 2.45 12.05 8.85 ;
        RECT  11.55 3.55 12.25 4.25 ;
        RECT  11.55 7.15 12.25 8.85 ;
    END
END NO4I3X1
MACRO NO4I3X2
    CLASS CORE ;
    FOREIGN NO4I3X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  14.25 2.55 14.75 10.50 ;
        RECT  14.25 7.10 14.95 10.50 ;
        RECT  14.25 2.55 15.15 4.20 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  9.55 5.40 10.95 6.15 ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  12.35 5.40 13.75 6.30 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 3.05 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.90 2.50 11.00 ;
        RECT  4.65 7.90 5.35 11.00 ;
        RECT  3.30 10.10 5.90 11.00 ;
        RECT  7.50 7.70 8.20 11.00 ;
        RECT  11.35 10.20 12.05 11.00 ;
        RECT  12.90 7.30 13.60 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.15 2.00 2.85 4.25 ;
        RECT  2.00 3.55 2.85 4.25 ;
        RECT  4.80 4.10 5.50 4.80 ;
        RECT  6.05 2.00 6.55 4.60 ;
        RECT  4.80 4.10 6.55 4.60 ;
        RECT  7.15 2.00 7.85 3.10 ;
        RECT  9.85 2.00 10.55 3.10 ;
        RECT  12.90 2.00 13.60 4.20 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.30 2.45 0.80 9.55 ;
        RECT  0.30 2.45 1.00 4.25 ;
        RECT  0.30 7.95 1.15 9.55 ;
        RECT  0.30 3.55 1.35 4.25 ;
        RECT  1.25 6.75 1.95 7.45 ;
        RECT  1.25 6.75 4.00 7.25 ;
        RECT  3.50 2.50 4.00 8.50 ;
        RECT  3.30 6.75 4.00 8.50 ;
        RECT  3.50 2.50 5.20 3.20 ;
        RECT  6.00 7.85 6.85 8.55 ;
        RECT  6.35 5.45 6.70 10.55 ;
        RECT  6.20 5.45 6.70 8.55 ;
        RECT  6.35 7.85 6.85 10.55 ;
        RECT  6.35 9.85 7.05 10.55 ;
        RECT  7.15 4.10 7.65 5.95 ;
        RECT  6.20 5.45 7.65 5.95 ;
        RECT  7.15 4.10 7.85 4.85 ;
        RECT  7.15 6.40 7.85 7.25 ;
        RECT  8.50 2.45 9.00 7.25 ;
        RECT  8.50 2.45 9.20 3.15 ;
        RECT  7.15 6.75 10.35 7.25 ;
        RECT  9.85 6.75 10.35 10.45 ;
        RECT  9.85 7.55 10.55 10.45 ;
        RECT  11.05 2.45 11.90 3.15 ;
        RECT  11.40 2.45 11.90 8.85 ;
        RECT  11.40 3.55 12.10 4.25 ;
        RECT  11.40 7.15 12.10 8.85 ;
    END
END NO4I3X2
MACRO NO4I3X4
    CLASS CORE ;
    FOREIGN NO4I3X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  14.25 2.55 14.75 10.50 ;
        RECT  14.25 7.10 14.95 10.50 ;
        RECT  14.25 2.55 15.15 4.20 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  9.55 5.40 10.95 6.15 ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  12.35 5.40 13.75 6.30 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 3.05 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.90 2.50 11.00 ;
        RECT  4.65 7.90 5.35 11.00 ;
        RECT  3.30 10.10 5.90 11.00 ;
        RECT  7.50 7.70 8.20 11.00 ;
        RECT  11.35 10.20 12.05 11.00 ;
        RECT  12.90 7.30 13.60 11.00 ;
        RECT  15.60 7.30 16.30 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.15 2.00 2.85 4.25 ;
        RECT  2.00 3.55 2.85 4.25 ;
        RECT  5.65 2.00 6.15 4.80 ;
        RECT  4.80 4.10 6.15 4.80 ;
        RECT  7.15 2.00 7.85 3.10 ;
        RECT  9.85 2.00 10.55 3.10 ;
        RECT  12.90 2.00 13.60 4.20 ;
        RECT  15.60 2.00 16.30 4.20 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.30 2.45 0.80 9.55 ;
        RECT  0.30 2.45 1.00 4.25 ;
        RECT  0.30 7.95 1.15 9.55 ;
        RECT  0.30 3.55 1.35 4.25 ;
        RECT  1.25 6.75 1.95 7.45 ;
        RECT  1.25 6.75 4.00 7.25 ;
        RECT  3.50 2.50 4.00 8.50 ;
        RECT  3.30 6.75 4.00 8.50 ;
        RECT  3.50 2.50 5.20 3.20 ;
        RECT  6.00 7.85 6.85 8.55 ;
        RECT  6.35 5.45 6.70 10.55 ;
        RECT  6.20 5.45 6.70 8.55 ;
        RECT  6.35 7.85 6.85 10.55 ;
        RECT  6.35 9.85 7.05 10.55 ;
        RECT  7.15 4.10 7.65 5.95 ;
        RECT  6.20 5.45 7.65 5.95 ;
        RECT  7.15 4.10 7.85 4.85 ;
        RECT  7.15 6.40 7.85 7.25 ;
        RECT  8.50 2.45 9.00 7.25 ;
        RECT  8.50 2.45 9.20 3.15 ;
        RECT  7.15 6.75 10.35 7.25 ;
        RECT  9.85 6.75 10.35 10.45 ;
        RECT  9.85 7.55 10.55 10.45 ;
        RECT  11.05 2.45 11.90 3.15 ;
        RECT  11.40 2.45 11.90 8.85 ;
        RECT  11.40 3.55 12.10 4.25 ;
        RECT  11.40 7.15 12.10 8.85 ;
    END
END NO4I3X4
MACRO NO4X1
    CLASS CORE ;
    FOREIGN NO4X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.45 2.60 11.95 9.15 ;
        RECT  10.30 8.45 11.95 9.15 ;
        RECT  11.45 2.60 12.35 3.70 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  9.55 3.85 10.95 4.55 ;
        RECT  10.05 3.85 10.95 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  8.30 5.40 9.55 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.45 2.55 7.60 ;
        RECT  1.65 6.45 2.90 7.15 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.00 7.65 3.70 11.00 ;
        RECT  5.85 7.55 6.55 11.00 ;
        RECT  9.35 7.30 9.85 10.30 ;
        RECT  9.35 9.80 10.90 10.30 ;
        RECT  10.20 7.10 10.90 7.80 ;
        RECT  9.35 7.30 10.90 7.80 ;
        RECT  10.05 9.80 10.90 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.20 ;
        RECT  3.20 2.50 4.15 3.20 ;
        RECT  3.55 2.00 4.15 4.80 ;
        RECT  3.45 4.10 4.15 4.80 ;
        RECT  4.85 2.00 6.45 2.90 ;
        RECT  7.40 2.00 8.10 3.20 ;
        RECT  10.10 2.00 10.80 3.25 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.55 5.45 1.05 10.05 ;
        RECT  0.45 7.55 1.15 10.05 ;
        RECT  1.60 2.55 2.10 5.95 ;
        RECT  1.60 2.55 2.50 3.25 ;
        RECT  0.55 5.45 4.10 5.95 ;
        RECT  3.40 5.35 4.10 6.05 ;
        RECT  4.50 7.55 5.20 8.25 ;
        RECT  4.70 4.35 5.10 10.15 ;
        RECT  4.60 4.35 5.10 8.25 ;
        RECT  4.70 7.55 5.20 10.15 ;
        RECT  4.70 9.45 5.40 10.15 ;
        RECT  5.55 5.35 6.25 6.05 ;
        RECT  5.80 4.10 6.50 4.85 ;
        RECT  4.60 4.35 6.50 4.85 ;
        RECT  5.55 5.35 7.85 5.85 ;
        RECT  7.35 3.75 7.85 8.05 ;
        RECT  7.35 7.55 8.90 8.05 ;
        RECT  8.20 7.55 8.90 10.05 ;
        RECT  8.60 2.50 9.10 4.25 ;
        RECT  7.35 3.75 9.10 4.25 ;
        RECT  8.60 2.50 9.50 3.30 ;
    END
END NO4X1
MACRO NO4X2
    CLASS CORE ;
    FOREIGN NO4X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.45 2.45 11.95 10.50 ;
        RECT  11.25 7.10 11.95 10.50 ;
        RECT  11.45 2.45 12.35 4.10 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  9.55 5.40 10.95 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  7.25 4.10 8.15 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.45 2.55 7.60 ;
        RECT  1.65 6.45 2.90 7.15 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.00 7.65 3.70 11.00 ;
        RECT  6.00 7.55 6.70 11.00 ;
        RECT  9.90 7.30 10.60 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.20 ;
        RECT  3.20 2.00 4.05 3.20 ;
        RECT  3.35 2.00 4.05 4.80 ;
        RECT  4.85 2.00 6.45 2.90 ;
        RECT  7.25 2.00 7.95 3.15 ;
        RECT  10.10 2.00 10.80 4.10 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.50 7.55 5.20 8.25 ;
        RECT  0.55 5.45 1.05 10.05 ;
        RECT  0.45 7.55 1.15 10.05 ;
        RECT  1.80 2.55 2.30 5.95 ;
        RECT  1.80 2.55 2.50 3.25 ;
        RECT  0.55 5.45 4.05 5.95 ;
        RECT  3.35 5.35 4.05 6.05 ;
        RECT  4.70 4.35 5.00 10.55 ;
        RECT  4.50 4.35 5.00 8.25 ;
        RECT  4.70 7.55 5.20 10.55 ;
        RECT  4.70 9.85 5.40 10.55 ;
        RECT  5.45 5.35 6.15 6.05 ;
        RECT  5.70 4.10 6.40 4.85 ;
        RECT  4.50 4.35 6.40 4.85 ;
        RECT  8.60 2.45 8.90 10.05 ;
        RECT  8.35 5.55 8.90 10.05 ;
        RECT  8.35 7.55 9.05 10.05 ;
        RECT  8.60 2.45 9.10 6.05 ;
        RECT  5.45 5.55 9.10 6.05 ;
        RECT  8.60 2.45 9.30 3.15 ;
    END
END NO4X2
MACRO NO4X3
    CLASS CORE ;
    FOREIGN NO4X3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.30 3.10 12.00 3.80 ;
        RECT  11.45 3.10 11.95 9.65 ;
        RECT  11.45 3.10 12.00 5.00 ;
        RECT  11.30 7.10 12.00 9.65 ;
        RECT  11.45 4.10 12.35 5.00 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  9.55 5.40 10.95 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  7.25 4.10 8.15 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.45 2.55 7.60 ;
        RECT  1.65 6.45 2.90 7.15 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.00 7.65 3.70 11.00 ;
        RECT  6.00 7.55 6.70 11.00 ;
        RECT  9.95 7.30 10.65 11.00 ;
        RECT  12.65 7.30 13.35 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.20 ;
        RECT  3.20 2.00 4.05 3.20 ;
        RECT  3.35 2.00 4.05 4.80 ;
        RECT  4.85 2.00 6.45 2.90 ;
        RECT  7.25 2.00 7.95 3.65 ;
        RECT  9.95 2.00 10.65 3.60 ;
        RECT  12.65 2.00 13.35 3.70 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.50 7.55 5.20 8.25 ;
        RECT  0.55 5.45 1.05 10.05 ;
        RECT  0.45 7.55 1.15 10.05 ;
        RECT  1.80 2.55 2.30 5.95 ;
        RECT  1.80 2.55 2.50 3.25 ;
        RECT  0.55 5.45 4.05 5.95 ;
        RECT  3.35 5.35 4.05 6.05 ;
        RECT  4.70 4.35 5.00 10.55 ;
        RECT  4.50 4.35 5.00 8.25 ;
        RECT  4.70 7.55 5.20 10.55 ;
        RECT  4.70 9.85 5.40 10.55 ;
        RECT  5.45 5.35 6.15 6.05 ;
        RECT  5.70 4.10 6.40 4.85 ;
        RECT  4.50 4.35 6.40 4.85 ;
        RECT  8.60 2.95 8.90 10.05 ;
        RECT  8.35 5.55 8.90 10.05 ;
        RECT  8.35 7.55 9.05 10.05 ;
        RECT  8.60 2.95 9.10 6.05 ;
        RECT  5.45 5.55 9.10 6.05 ;
        RECT  8.60 2.95 9.30 3.65 ;
    END
END NO4X3
MACRO NO4X4
    CLASS CORE ;
    FOREIGN NO4X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.45 2.55 11.95 10.55 ;
        RECT  11.30 7.10 12.00 10.55 ;
        RECT  11.45 2.55 12.15 5.00 ;
        RECT  11.45 4.10 12.35 5.00 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  9.55 5.40 10.95 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  7.25 4.10 8.15 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.45 2.55 7.60 ;
        RECT  1.65 6.45 2.90 7.15 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.00 7.65 3.70 11.00 ;
        RECT  6.00 7.55 6.70 11.00 ;
        RECT  9.95 7.30 10.65 11.00 ;
        RECT  12.65 7.30 13.35 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.20 ;
        RECT  3.20 2.00 4.05 3.20 ;
        RECT  3.35 2.00 4.05 4.80 ;
        RECT  4.85 2.00 6.45 2.90 ;
        RECT  7.25 2.00 7.95 3.65 ;
        RECT  10.10 2.00 10.80 4.15 ;
        RECT  12.80 2.00 13.50 4.15 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.50 7.55 5.20 8.25 ;
        RECT  0.55 5.45 1.05 10.05 ;
        RECT  0.45 7.55 1.15 10.05 ;
        RECT  1.80 2.55 2.30 5.95 ;
        RECT  1.80 2.55 2.50 3.25 ;
        RECT  0.55 5.45 4.05 5.95 ;
        RECT  3.35 5.35 4.05 6.05 ;
        RECT  4.70 4.35 5.00 10.55 ;
        RECT  4.50 4.35 5.00 8.25 ;
        RECT  4.70 7.55 5.20 10.55 ;
        RECT  4.70 9.85 5.40 10.55 ;
        RECT  5.45 5.35 6.15 6.05 ;
        RECT  5.70 4.10 6.40 4.85 ;
        RECT  4.50 4.35 6.40 4.85 ;
        RECT  8.60 2.95 8.90 10.05 ;
        RECT  8.35 5.55 8.90 10.05 ;
        RECT  8.35 7.55 9.05 10.05 ;
        RECT  8.60 2.95 9.10 6.05 ;
        RECT  5.45 5.55 9.10 6.05 ;
        RECT  8.60 2.95 9.30 3.65 ;
    END
END NO4X4
MACRO NO5I1X1
    CLASS CORE ;
    FOREIGN NO5I1X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  15.65 2.80 16.15 8.75 ;
        RECT  15.65 7.15 16.35 8.75 ;
        RECT  15.65 2.80 16.55 3.70 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  13.85 5.40 15.15 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  11.45 4.10 12.35 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  5.65 5.30 6.75 6.00 ;
        RECT  5.85 5.30 6.75 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.45 4.65 3.95 6.30 ;
        RECT  3.05 5.40 3.95 6.30 ;
        RECT  3.45 4.65 4.25 5.35 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 10.10 1.15 11.00 ;
        RECT  1.95 7.70 2.65 11.00 ;
        RECT  6.80 7.70 7.50 11.00 ;
        RECT  9.65 7.20 10.35 11.00 ;
        RECT  14.25 7.30 14.95 11.00 ;
        RECT  13.75 10.10 16.35 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 3.25 ;
        RECT  4.50 2.00 5.20 3.25 ;
        RECT  7.35 2.00 8.05 3.65 ;
        RECT  11.60 2.00 12.30 3.65 ;
        RECT  14.30 2.00 15.00 3.65 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 2.60 1.15 3.30 ;
        RECT  0.65 2.60 1.15 4.20 ;
        RECT  0.45 6.75 1.15 9.10 ;
        RECT  0.65 3.70 2.15 4.20 ;
        RECT  1.65 3.70 2.15 7.25 ;
        RECT  0.45 6.75 2.15 7.25 ;
        RECT  1.65 5.30 2.60 6.00 ;
        RECT  3.15 2.60 3.85 4.20 ;
        RECT  4.70 3.70 5.20 7.25 ;
        RECT  5.30 6.75 6.00 10.55 ;
        RECT  5.85 2.60 6.55 4.20 ;
        RECT  3.15 3.70 6.55 4.20 ;
        RECT  7.20 6.55 7.90 7.25 ;
        RECT  4.70 6.75 7.90 7.25 ;
        RECT  8.15 7.70 8.85 8.40 ;
        RECT  8.35 4.45 8.85 10.55 ;
        RECT  8.35 9.85 9.20 10.55 ;
        RECT  9.30 5.45 10.00 6.15 ;
        RECT  9.70 3.00 10.20 5.00 ;
        RECT  8.35 4.45 10.20 5.00 ;
        RECT  9.70 3.00 10.40 3.70 ;
        RECT  12.00 5.45 12.50 10.55 ;
        RECT  12.00 7.15 12.70 10.55 ;
        RECT  12.80 3.00 13.30 5.95 ;
        RECT  9.30 5.45 13.30 5.95 ;
        RECT  12.80 3.00 13.65 3.70 ;
    END
END NO5I1X1
MACRO NO5I1X2
    CLASS CORE ;
    FOREIGN NO5I1X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  15.65 2.75 16.15 10.55 ;
        RECT  15.65 7.15 16.35 10.55 ;
        RECT  15.65 2.75 16.55 4.40 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  13.85 5.40 15.15 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  11.45 4.10 12.35 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  5.65 5.30 6.75 6.00 ;
        RECT  5.85 5.30 6.75 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.45 4.65 3.95 6.30 ;
        RECT  3.05 5.40 3.95 6.30 ;
        RECT  3.45 4.65 4.25 5.35 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 10.10 1.15 11.00 ;
        RECT  1.95 7.70 2.65 11.00 ;
        RECT  6.80 7.70 7.50 11.00 ;
        RECT  9.65 7.20 10.35 11.00 ;
        RECT  14.25 7.30 14.95 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 3.25 ;
        RECT  4.50 2.00 5.20 3.25 ;
        RECT  7.35 2.00 8.05 3.65 ;
        RECT  11.45 2.00 12.15 3.65 ;
        RECT  14.30 2.00 15.00 4.40 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 2.60 1.15 3.30 ;
        RECT  0.65 2.60 1.15 4.20 ;
        RECT  0.45 6.75 1.15 9.10 ;
        RECT  0.65 3.70 2.15 4.20 ;
        RECT  1.65 3.70 2.15 7.25 ;
        RECT  0.45 6.75 2.15 7.25 ;
        RECT  1.65 5.30 2.60 6.00 ;
        RECT  3.15 2.60 3.85 4.20 ;
        RECT  4.70 3.70 5.20 7.25 ;
        RECT  5.30 6.75 6.00 10.55 ;
        RECT  5.85 2.60 6.55 4.20 ;
        RECT  3.15 3.70 6.55 4.20 ;
        RECT  7.20 6.55 7.90 7.25 ;
        RECT  4.70 6.75 7.90 7.25 ;
        RECT  8.15 7.70 8.85 8.40 ;
        RECT  8.35 4.45 8.85 10.55 ;
        RECT  8.35 9.85 9.20 10.55 ;
        RECT  9.30 5.45 10.00 6.15 ;
        RECT  9.70 3.00 10.20 5.00 ;
        RECT  8.35 4.45 10.20 5.00 ;
        RECT  9.70 3.00 10.40 3.70 ;
        RECT  12.00 5.45 12.50 10.55 ;
        RECT  12.00 7.15 12.70 10.55 ;
        RECT  12.80 3.00 13.30 5.95 ;
        RECT  9.30 5.45 13.30 5.95 ;
        RECT  12.80 3.00 13.50 3.70 ;
    END
END NO5I1X2
MACRO NO5I1X4
    CLASS CORE ;
    FOREIGN NO5I1X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  15.65 2.75 16.15 10.55 ;
        RECT  15.65 7.15 16.35 10.55 ;
        RECT  15.65 2.75 16.55 4.40 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  13.85 5.40 15.15 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  11.45 4.10 12.35 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  5.65 5.30 6.75 6.00 ;
        RECT  5.85 5.30 6.75 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.45 4.65 3.95 6.30 ;
        RECT  3.05 5.40 3.95 6.30 ;
        RECT  3.45 4.65 4.25 5.35 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 10.10 1.15 11.00 ;
        RECT  1.95 7.70 2.65 11.00 ;
        RECT  6.80 7.70 7.50 11.00 ;
        RECT  9.65 7.20 10.35 11.00 ;
        RECT  14.30 7.30 15.00 11.00 ;
        RECT  17.00 7.30 17.70 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 3.25 ;
        RECT  4.50 2.00 5.20 3.25 ;
        RECT  7.35 2.00 8.05 3.65 ;
        RECT  11.45 2.00 12.15 3.65 ;
        RECT  14.30 2.00 15.00 4.40 ;
        RECT  17.00 2.00 17.70 4.40 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 2.60 1.15 3.30 ;
        RECT  0.65 2.60 1.15 4.20 ;
        RECT  0.45 6.75 1.15 9.10 ;
        RECT  0.65 3.70 2.15 4.20 ;
        RECT  1.65 3.70 2.15 7.25 ;
        RECT  0.45 6.75 2.15 7.25 ;
        RECT  1.65 5.30 2.60 6.00 ;
        RECT  3.15 2.60 3.85 4.20 ;
        RECT  4.70 3.70 5.20 7.25 ;
        RECT  5.30 6.75 6.00 10.55 ;
        RECT  5.85 2.60 6.55 4.20 ;
        RECT  3.15 3.70 6.55 4.20 ;
        RECT  7.20 6.55 7.90 7.25 ;
        RECT  4.70 6.75 7.90 7.25 ;
        RECT  8.15 7.70 8.85 8.40 ;
        RECT  8.35 4.45 8.85 10.55 ;
        RECT  8.35 9.85 9.20 10.55 ;
        RECT  9.30 5.45 10.00 6.15 ;
        RECT  9.70 3.00 10.20 5.00 ;
        RECT  8.35 4.45 10.20 5.00 ;
        RECT  9.70 3.00 10.40 3.70 ;
        RECT  12.00 5.45 12.50 10.55 ;
        RECT  12.00 7.15 12.70 10.55 ;
        RECT  12.80 3.00 13.30 5.95 ;
        RECT  9.30 5.45 13.30 5.95 ;
        RECT  12.80 3.00 13.50 3.70 ;
    END
END NO5I1X4
MACRO NO5I2X1
    CLASS CORE ;
    FOREIGN NO5I2X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  15.65 2.45 16.00 8.80 ;
        RECT  15.30 2.45 16.00 3.70 ;
        RECT  15.65 2.80 16.15 8.80 ;
        RECT  15.65 7.20 16.35 8.80 ;
        RECT  15.30 2.80 16.55 3.70 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  13.75 5.40 15.15 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  10.30 4.65 11.00 6.30 ;
        RECT  10.05 5.40 11.00 6.30 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 3.05 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.90 2.50 11.00 ;
        RECT  4.65 7.90 5.35 11.00 ;
        RECT  3.30 10.10 6.70 11.00 ;
        RECT  7.65 7.80 8.35 11.00 ;
        RECT  14.30 7.20 15.00 11.00 ;
        RECT  14.30 10.10 16.35 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.00 2.00 2.70 4.45 ;
        RECT  5.85 2.00 6.55 4.45 ;
        RECT  11.25 2.00 11.95 3.15 ;
        RECT  13.95 2.00 14.65 3.20 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 2.45 0.95 9.55 ;
        RECT  0.30 2.45 1.00 3.15 ;
        RECT  0.45 7.95 1.15 9.55 ;
        RECT  0.45 3.75 1.35 4.45 ;
        RECT  1.40 6.75 2.10 7.45 ;
        RECT  1.40 6.75 4.00 7.25 ;
        RECT  3.50 3.70 4.00 8.50 ;
        RECT  3.30 6.75 4.00 8.50 ;
        RECT  3.50 3.70 5.05 4.40 ;
        RECT  6.15 5.60 6.65 8.55 ;
        RECT  6.15 7.85 6.85 8.55 ;
        RECT  7.20 6.55 7.90 7.25 ;
        RECT  8.20 3.75 8.70 6.10 ;
        RECT  8.40 2.45 8.70 6.10 ;
        RECT  6.15 5.60 8.70 6.10 ;
        RECT  8.40 2.45 8.90 4.45 ;
        RECT  8.20 3.75 8.90 4.45 ;
        RECT  8.40 2.45 9.25 3.15 ;
        RECT  9.90 2.45 10.60 3.15 ;
        RECT  10.10 2.45 10.60 4.10 ;
        RECT  12.60 2.45 13.30 3.15 ;
        RECT  10.10 3.60 13.30 4.10 ;
        RECT  7.20 6.75 13.30 7.25 ;
        RECT  11.00 8.20 13.50 8.90 ;
        RECT  12.80 2.45 13.30 10.50 ;
        RECT  12.80 8.20 13.50 10.50 ;
    END
END NO5I2X1
MACRO NO5I2X2
    CLASS CORE ;
    FOREIGN NO5I2X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  15.65 2.45 16.15 10.50 ;
        RECT  15.65 7.10 16.35 10.50 ;
        RECT  15.50 2.45 16.55 4.10 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  13.75 5.40 15.15 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  10.30 4.65 11.00 6.30 ;
        RECT  10.05 5.40 11.00 6.30 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 3.05 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.90 2.50 11.00 ;
        RECT  4.65 7.90 5.35 11.00 ;
        RECT  3.30 10.10 6.70 11.00 ;
        RECT  7.65 7.80 8.35 11.00 ;
        RECT  14.30 7.30 15.00 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.00 2.00 2.70 4.45 ;
        RECT  5.85 2.00 6.55 4.45 ;
        RECT  11.25 2.00 11.95 3.15 ;
        RECT  14.15 2.00 14.85 4.10 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 2.45 0.95 9.55 ;
        RECT  0.30 2.45 1.00 3.15 ;
        RECT  0.45 7.95 1.15 9.55 ;
        RECT  0.45 3.75 1.35 4.45 ;
        RECT  1.40 6.75 2.10 7.45 ;
        RECT  1.40 6.75 4.00 7.25 ;
        RECT  3.50 3.70 4.00 8.50 ;
        RECT  3.30 6.75 4.00 8.50 ;
        RECT  3.50 3.70 5.05 4.40 ;
        RECT  6.15 5.60 6.65 8.55 ;
        RECT  6.15 7.85 6.85 8.55 ;
        RECT  7.20 6.55 7.90 7.25 ;
        RECT  8.20 3.75 8.70 6.10 ;
        RECT  8.40 2.45 8.70 6.10 ;
        RECT  6.15 5.60 8.70 6.10 ;
        RECT  8.40 2.45 8.90 4.45 ;
        RECT  8.20 3.75 8.90 4.45 ;
        RECT  8.40 2.45 9.25 3.15 ;
        RECT  9.90 2.45 10.60 3.15 ;
        RECT  10.10 2.45 10.60 4.10 ;
        RECT  12.60 2.45 13.30 3.15 ;
        RECT  10.10 3.60 13.30 4.10 ;
        RECT  7.20 6.75 13.30 7.25 ;
        RECT  11.00 8.20 13.50 8.90 ;
        RECT  12.80 2.45 13.30 10.50 ;
        RECT  12.80 8.20 13.50 10.50 ;
    END
END NO5I2X2
MACRO NO5I2X4
    CLASS CORE ;
    FOREIGN NO5I2X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  15.65 2.45 16.15 10.50 ;
        RECT  15.50 2.45 16.20 4.10 ;
        RECT  15.65 7.10 16.35 10.50 ;
        RECT  15.65 8.00 16.55 8.90 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  13.75 5.40 15.15 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  10.30 4.65 11.00 6.30 ;
        RECT  10.05 5.40 11.00 6.30 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 3.05 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.90 2.50 11.00 ;
        RECT  4.65 7.90 5.35 11.00 ;
        RECT  3.30 10.10 6.70 11.00 ;
        RECT  7.65 7.80 8.35 11.00 ;
        RECT  14.30 7.30 15.00 11.00 ;
        RECT  17.00 7.30 17.70 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.00 2.00 2.70 4.45 ;
        RECT  5.85 2.00 6.55 4.45 ;
        RECT  11.25 2.00 11.95 3.15 ;
        RECT  14.15 2.00 14.85 4.10 ;
        RECT  16.85 2.00 17.55 4.10 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 2.45 0.95 9.55 ;
        RECT  0.30 2.45 1.00 3.15 ;
        RECT  0.45 7.95 1.15 9.55 ;
        RECT  0.45 3.75 1.35 4.45 ;
        RECT  1.40 6.75 2.10 7.45 ;
        RECT  1.40 6.75 4.00 7.25 ;
        RECT  3.50 3.70 4.00 8.50 ;
        RECT  3.30 6.75 4.00 8.50 ;
        RECT  3.50 3.70 5.05 4.40 ;
        RECT  6.15 5.60 6.65 8.55 ;
        RECT  6.15 7.85 6.85 8.55 ;
        RECT  7.20 6.55 7.90 7.25 ;
        RECT  8.20 3.75 8.70 6.10 ;
        RECT  8.40 2.45 8.70 6.10 ;
        RECT  6.15 5.60 8.70 6.10 ;
        RECT  8.40 2.45 8.90 4.45 ;
        RECT  8.20 3.75 8.90 4.45 ;
        RECT  8.40 2.45 9.25 3.15 ;
        RECT  9.90 2.45 10.60 3.15 ;
        RECT  10.10 2.45 10.60 4.10 ;
        RECT  12.60 2.45 13.30 3.15 ;
        RECT  10.10 3.60 13.30 4.10 ;
        RECT  7.20 6.75 13.30 7.25 ;
        RECT  11.00 8.20 13.50 8.90 ;
        RECT  12.80 2.45 13.30 10.50 ;
        RECT  12.80 8.20 13.50 10.50 ;
    END
END NO5I2X4
MACRO NO5I3X1
    CLASS CORE ;
    FOREIGN NO5I3X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  14.25 2.80 14.75 8.80 ;
        RECT  14.25 7.10 14.95 8.80 ;
        RECT  14.25 2.80 15.15 3.70 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  12.45 5.40 13.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  10.05 4.10 10.95 5.00 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 4.40 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.55 7.60 ;
        RECT  1.65 6.75 2.90 7.60 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.05 2.50 11.00 ;
        RECT  3.50 7.50 4.20 11.00 ;
        RECT  6.20 7.55 6.90 11.00 ;
        RECT  6.20 10.10 7.45 11.00 ;
        RECT  9.05 7.55 9.75 11.00 ;
        RECT  12.90 7.15 13.60 11.00 ;
        RECT  12.90 10.10 14.95 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.70 2.00 3.40 3.20 ;
        RECT  6.20 4.05 6.90 4.75 ;
        RECT  7.40 2.00 7.90 4.55 ;
        RECT  6.20 4.05 7.90 4.55 ;
        RECT  7.40 2.00 9.40 2.90 ;
        RECT  10.20 2.00 10.90 3.65 ;
        RECT  12.90 2.00 13.60 3.65 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.30 2.45 0.80 9.70 ;
        RECT  0.30 8.10 1.15 9.70 ;
        RECT  0.30 2.45 2.05 3.15 ;
        RECT  1.35 3.70 2.05 4.40 ;
        RECT  1.35 3.70 5.35 4.20 ;
        RECT  4.85 2.70 5.35 10.55 ;
        RECT  4.85 7.50 5.55 8.20 ;
        RECT  4.85 9.85 5.55 10.55 ;
        RECT  6.05 2.50 6.75 3.20 ;
        RECT  4.85 2.70 6.75 3.20 ;
        RECT  7.55 7.55 8.40 8.25 ;
        RECT  7.90 5.45 8.15 10.55 ;
        RECT  7.65 5.45 8.15 8.25 ;
        RECT  7.90 7.55 8.40 10.55 ;
        RECT  7.90 9.85 8.60 10.55 ;
        RECT  8.55 4.05 9.05 5.95 ;
        RECT  7.65 5.45 9.05 5.95 ;
        RECT  8.55 4.05 9.25 4.80 ;
        RECT  8.60 6.40 9.30 7.10 ;
        RECT  8.60 6.60 11.90 7.10 ;
        RECT  11.40 2.95 11.90 10.45 ;
        RECT  11.40 7.55 12.10 10.45 ;
        RECT  11.40 2.95 12.25 3.65 ;
    END
END NO5I3X1
MACRO NO5I3X2
    CLASS CORE ;
    FOREIGN NO5I3X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  14.25 2.45 14.75 10.50 ;
        RECT  14.25 7.10 14.95 10.50 ;
        RECT  14.25 2.45 15.15 4.10 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  12.35 5.40 13.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  10.05 4.10 10.95 5.00 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 4.40 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.55 7.60 ;
        RECT  1.65 6.75 2.90 7.60 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.05 2.50 11.00 ;
        RECT  3.50 7.50 4.20 11.00 ;
        RECT  6.20 7.55 6.90 11.00 ;
        RECT  6.20 10.10 7.45 11.00 ;
        RECT  9.05 7.55 9.75 11.00 ;
        RECT  12.90 7.30 13.60 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.70 2.00 3.40 3.20 ;
        RECT  6.20 4.05 6.90 4.75 ;
        RECT  7.40 2.00 7.90 4.55 ;
        RECT  6.20 4.05 7.90 4.55 ;
        RECT  7.40 2.00 8.50 2.90 ;
        RECT  10.05 2.00 10.75 3.65 ;
        RECT  12.90 2.00 13.60 4.10 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.30 2.45 0.80 9.70 ;
        RECT  0.30 8.10 1.15 9.70 ;
        RECT  0.30 2.45 2.05 3.15 ;
        RECT  1.35 3.70 2.05 4.40 ;
        RECT  1.35 3.70 5.35 4.20 ;
        RECT  4.85 2.70 5.35 10.55 ;
        RECT  4.85 7.50 5.55 8.20 ;
        RECT  4.85 9.85 5.55 10.55 ;
        RECT  6.05 2.50 6.75 3.20 ;
        RECT  4.85 2.70 6.75 3.20 ;
        RECT  7.55 7.55 8.40 8.25 ;
        RECT  7.90 5.45 8.15 10.55 ;
        RECT  7.65 5.45 8.15 8.25 ;
        RECT  7.90 7.55 8.40 10.55 ;
        RECT  7.90 9.85 8.60 10.55 ;
        RECT  8.55 4.05 9.05 5.95 ;
        RECT  7.65 5.45 9.05 5.95 ;
        RECT  8.55 4.05 9.25 4.80 ;
        RECT  8.60 6.40 9.30 7.10 ;
        RECT  8.60 6.60 11.90 7.10 ;
        RECT  11.40 2.95 11.90 10.45 ;
        RECT  11.40 2.95 12.10 3.65 ;
        RECT  11.40 7.55 12.10 10.45 ;
    END
END NO5I3X2
MACRO NO5I3X4
    CLASS CORE ;
    FOREIGN NO5I3X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  14.25 2.75 14.75 10.50 ;
        RECT  14.25 7.10 14.95 10.50 ;
        RECT  14.25 2.75 15.15 4.40 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  12.35 5.40 13.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  10.05 4.10 10.95 5.00 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 4.40 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.55 7.60 ;
        RECT  1.65 6.75 2.90 7.60 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.05 2.50 11.00 ;
        RECT  3.50 7.50 4.20 11.00 ;
        RECT  6.20 7.55 6.90 11.00 ;
        RECT  6.20 10.10 7.45 11.00 ;
        RECT  9.05 7.55 9.75 11.00 ;
        RECT  12.90 7.30 13.60 11.00 ;
        RECT  15.60 7.30 16.30 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.70 2.00 3.40 3.20 ;
        RECT  6.20 4.05 6.90 4.75 ;
        RECT  7.40 2.00 7.90 4.55 ;
        RECT  6.20 4.05 7.90 4.55 ;
        RECT  7.40 2.00 8.50 2.90 ;
        RECT  10.05 2.00 10.75 3.65 ;
        RECT  12.90 2.00 13.60 4.40 ;
        RECT  15.60 2.00 16.30 4.40 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.30 2.45 0.80 9.70 ;
        RECT  0.30 8.10 1.15 9.70 ;
        RECT  0.30 2.45 2.05 3.15 ;
        RECT  1.35 3.70 2.05 4.40 ;
        RECT  1.35 3.70 5.35 4.20 ;
        RECT  4.85 2.70 5.35 10.55 ;
        RECT  4.85 7.50 5.55 8.20 ;
        RECT  4.85 9.85 5.55 10.55 ;
        RECT  6.05 2.50 6.75 3.20 ;
        RECT  4.85 2.70 6.75 3.20 ;
        RECT  7.55 7.55 8.40 8.25 ;
        RECT  7.90 5.45 8.15 10.55 ;
        RECT  7.65 5.45 8.15 8.25 ;
        RECT  7.90 7.55 8.40 10.55 ;
        RECT  7.90 9.85 8.60 10.55 ;
        RECT  8.55 4.05 9.05 5.95 ;
        RECT  7.65 5.45 9.05 5.95 ;
        RECT  8.55 4.05 9.25 4.80 ;
        RECT  8.60 6.40 9.30 7.10 ;
        RECT  8.60 6.60 11.90 7.10 ;
        RECT  11.40 2.95 11.90 10.45 ;
        RECT  11.40 2.95 12.10 3.65 ;
        RECT  11.40 7.55 12.10 10.45 ;
    END
END NO5I3X4
MACRO NO5I4X1
    CLASS CORE ;
    FOREIGN NO5I4X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  15.65 2.80 16.15 8.80 ;
        RECT  15.65 7.20 16.35 8.80 ;
        RECT  15.65 2.80 16.55 4.25 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  11.45 4.10 12.35 5.00 ;
        END
    END E
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  13.95 5.40 15.15 6.30 ;
        END
    END DN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 4.40 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.55 7.60 ;
        RECT  1.65 6.75 2.90 7.60 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.05 2.50 11.00 ;
        RECT  3.50 7.50 4.20 11.00 ;
        RECT  6.20 7.55 6.90 11.00 ;
        RECT  6.20 10.10 7.45 11.00 ;
        RECT  9.05 7.55 9.75 11.00 ;
        RECT  14.30 7.20 15.00 11.00 ;
        RECT  13.20 10.50 16.25 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.70 2.00 3.40 3.20 ;
        RECT  6.20 4.05 6.90 4.75 ;
        RECT  7.40 2.00 7.90 4.55 ;
        RECT  6.20 4.05 7.90 4.55 ;
        RECT  8.60 2.00 9.30 3.10 ;
        RECT  11.30 2.00 12.00 3.10 ;
        RECT  14.30 2.00 15.00 4.25 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.30 2.45 0.80 9.70 ;
        RECT  0.30 8.10 1.15 9.70 ;
        RECT  0.30 2.45 2.05 3.15 ;
        RECT  1.35 3.70 2.05 4.40 ;
        RECT  1.35 3.70 5.35 4.20 ;
        RECT  4.85 2.70 5.35 10.55 ;
        RECT  4.85 7.50 5.55 8.20 ;
        RECT  4.85 9.85 5.55 10.55 ;
        RECT  6.05 2.50 6.75 3.20 ;
        RECT  4.85 2.70 6.75 3.20 ;
        RECT  7.55 7.55 8.40 8.25 ;
        RECT  7.90 5.45 8.15 10.55 ;
        RECT  7.65 5.45 8.15 8.25 ;
        RECT  7.90 7.55 8.40 10.55 ;
        RECT  7.90 9.85 8.60 10.55 ;
        RECT  8.55 4.10 9.05 5.95 ;
        RECT  7.65 5.45 9.05 5.95 ;
        RECT  8.55 4.10 9.25 4.80 ;
        RECT  8.60 6.40 9.30 7.10 ;
        RECT  9.95 2.45 10.65 3.15 ;
        RECT  10.15 2.45 10.65 7.10 ;
        RECT  8.60 6.60 11.90 7.10 ;
        RECT  11.40 6.60 11.90 10.45 ;
        RECT  11.40 7.55 12.10 10.45 ;
        RECT  12.45 2.45 13.45 3.15 ;
        RECT  12.95 2.45 13.45 8.80 ;
        RECT  12.95 3.55 13.65 4.25 ;
        RECT  12.95 7.20 13.65 8.80 ;
    END
END NO5I4X1
MACRO NO5I4X2
    CLASS CORE ;
    FOREIGN NO5I4X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  15.65 2.55 16.15 10.50 ;
        RECT  15.65 7.10 16.35 10.50 ;
        RECT  15.65 2.55 16.55 4.20 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  11.45 4.10 12.35 5.00 ;
        END
    END E
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  13.95 5.40 15.15 6.30 ;
        END
    END DN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 4.40 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.55 7.60 ;
        RECT  1.65 6.75 2.90 7.60 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.05 2.50 11.00 ;
        RECT  3.50 7.50 4.20 11.00 ;
        RECT  6.20 7.55 6.90 11.00 ;
        RECT  6.20 10.10 7.35 11.00 ;
        RECT  8.95 7.55 9.65 11.00 ;
        RECT  14.30 7.30 15.00 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.70 2.00 3.40 3.20 ;
        RECT  6.20 4.05 6.90 4.75 ;
        RECT  7.40 2.00 7.90 4.55 ;
        RECT  6.20 4.05 7.90 4.55 ;
        RECT  8.60 2.00 9.30 3.10 ;
        RECT  11.30 2.00 12.00 3.10 ;
        RECT  14.30 2.00 15.00 4.20 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.30 2.45 0.80 9.70 ;
        RECT  0.30 8.10 1.15 9.70 ;
        RECT  0.30 2.45 2.05 3.15 ;
        RECT  1.35 3.70 2.05 4.40 ;
        RECT  1.35 3.70 5.35 4.20 ;
        RECT  4.85 2.70 5.35 10.55 ;
        RECT  4.85 7.50 5.55 8.20 ;
        RECT  4.85 9.85 5.55 10.55 ;
        RECT  6.05 2.50 6.75 3.20 ;
        RECT  4.85 2.70 6.75 3.20 ;
        RECT  7.55 7.55 8.30 8.25 ;
        RECT  7.80 5.45 8.15 10.55 ;
        RECT  7.65 5.45 8.15 8.25 ;
        RECT  7.80 7.55 8.30 10.55 ;
        RECT  7.80 9.85 8.50 10.55 ;
        RECT  8.55 4.10 9.05 5.95 ;
        RECT  7.65 5.45 9.05 5.95 ;
        RECT  8.55 4.10 9.25 4.80 ;
        RECT  8.60 6.40 9.30 7.10 ;
        RECT  9.95 2.45 10.65 3.15 ;
        RECT  10.15 2.45 10.65 7.10 ;
        RECT  8.60 6.60 11.80 7.10 ;
        RECT  11.30 6.60 11.80 10.45 ;
        RECT  11.30 7.55 12.00 10.45 ;
        RECT  12.45 2.45 13.30 3.15 ;
        RECT  12.80 2.45 13.30 8.80 ;
        RECT  12.80 3.50 13.50 4.20 ;
        RECT  12.80 7.20 13.50 8.80 ;
    END
END NO5I4X2
MACRO NO5I4X4
    CLASS CORE ;
    FOREIGN NO5I4X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  15.65 2.55 16.15 10.50 ;
        RECT  15.65 7.10 16.35 10.50 ;
        RECT  15.65 2.55 16.55 4.20 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  11.45 4.10 12.35 5.00 ;
        END
    END E
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  13.95 5.40 15.15 6.30 ;
        END
    END DN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 4.40 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.55 7.60 ;
        RECT  1.65 6.75 2.90 7.60 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.05 2.50 11.00 ;
        RECT  3.50 7.50 4.20 11.00 ;
        RECT  6.20 7.55 6.90 11.00 ;
        RECT  6.20 10.10 7.35 11.00 ;
        RECT  8.95 7.55 9.65 11.00 ;
        RECT  14.30 7.30 15.00 11.00 ;
        RECT  17.00 7.30 17.70 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.70 2.00 3.40 3.20 ;
        RECT  6.20 4.05 6.90 4.75 ;
        RECT  7.40 2.00 7.90 4.55 ;
        RECT  6.20 4.05 7.90 4.55 ;
        RECT  8.60 2.00 9.30 3.10 ;
        RECT  11.30 2.00 12.00 3.10 ;
        RECT  14.30 2.00 15.00 4.20 ;
        RECT  17.00 2.00 17.70 4.20 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.30 2.45 0.80 9.70 ;
        RECT  0.30 8.10 1.15 9.70 ;
        RECT  0.30 2.45 2.05 3.15 ;
        RECT  1.35 3.70 2.05 4.40 ;
        RECT  1.35 3.70 5.35 4.20 ;
        RECT  4.85 2.70 5.35 10.55 ;
        RECT  4.85 7.50 5.55 8.20 ;
        RECT  4.85 9.85 5.55 10.55 ;
        RECT  6.05 2.50 6.75 3.20 ;
        RECT  4.85 2.70 6.75 3.20 ;
        RECT  7.55 7.55 8.30 8.25 ;
        RECT  7.80 5.45 8.15 10.55 ;
        RECT  7.65 5.45 8.15 8.25 ;
        RECT  7.80 7.55 8.30 10.55 ;
        RECT  7.80 9.85 8.50 10.55 ;
        RECT  8.55 4.10 9.05 5.95 ;
        RECT  7.65 5.45 9.05 5.95 ;
        RECT  8.55 4.10 9.25 4.80 ;
        RECT  8.60 6.40 9.30 7.10 ;
        RECT  9.95 2.45 10.65 3.15 ;
        RECT  10.15 2.45 10.65 7.10 ;
        RECT  8.60 6.60 11.80 7.10 ;
        RECT  11.30 6.60 11.80 10.45 ;
        RECT  11.30 7.55 12.00 10.45 ;
        RECT  12.45 2.45 13.30 3.15 ;
        RECT  12.80 2.45 13.30 8.80 ;
        RECT  12.80 3.50 13.50 4.20 ;
        RECT  12.80 7.20 13.50 8.80 ;
    END
END NO5I4X4
MACRO NO5X1
    CLASS CORE ;
    FOREIGN NO5X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  12.70 8.70 13.40 9.40 ;
        RECT  14.20 2.75 14.70 9.25 ;
        RECT  12.70 8.70 14.70 9.25 ;
        RECT  14.20 2.75 15.15 3.70 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  12.45 4.10 13.75 4.90 ;
        RECT  12.85 4.10 13.75 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  11.15 5.40 12.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.40 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 3.95 5.00 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  1.65 9.30 2.55 10.20 ;
        RECT  3.55 6.55 4.05 9.80 ;
        RECT  1.65 9.30 4.05 9.80 ;
        RECT  5.05 6.35 5.75 7.05 ;
        RECT  3.55 6.55 5.75 7.05 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  5.25 7.70 5.95 11.00 ;
        RECT  8.25 7.55 8.95 11.00 ;
        RECT  11.75 7.50 12.25 11.00 ;
        RECT  12.60 7.35 13.30 8.05 ;
        RECT  11.75 7.50 13.30 8.05 ;
        RECT  12.70 10.05 13.40 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.90 2.00 3.60 3.60 ;
        RECT  5.60 2.00 6.30 3.60 ;
        RECT  10.20 2.00 10.90 3.60 ;
        RECT  12.90 2.00 13.60 3.60 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  10.15 7.55 11.30 8.05 ;
        RECT  0.65 7.40 1.15 9.90 ;
        RECT  0.45 8.30 1.15 9.90 ;
        RECT  1.55 3.00 2.25 3.70 ;
        RECT  1.75 3.00 2.25 8.10 ;
        RECT  0.65 7.40 2.60 8.10 ;
        RECT  4.25 2.95 4.95 3.65 ;
        RECT  4.45 2.95 4.70 5.95 ;
        RECT  1.75 5.45 4.70 5.95 ;
        RECT  4.45 2.95 4.95 5.90 ;
        RECT  1.75 5.45 4.95 5.90 ;
        RECT  4.45 5.25 6.75 5.75 ;
        RECT  6.05 5.05 6.75 5.75 ;
        RECT  1.75 5.45 6.75 5.75 ;
        RECT  6.75 7.55 7.75 8.25 ;
        RECT  7.25 3.10 7.75 10.55 ;
        RECT  7.05 9.85 7.75 10.55 ;
        RECT  7.95 2.95 8.65 3.65 ;
        RECT  7.25 3.10 8.65 3.65 ;
        RECT  8.30 4.20 9.00 4.90 ;
        RECT  10.60 4.20 10.65 10.05 ;
        RECT  10.15 4.20 10.65 8.05 ;
        RECT  10.60 7.55 11.30 10.05 ;
        RECT  11.50 2.95 12.00 4.70 ;
        RECT  8.30 4.20 12.00 4.70 ;
        RECT  11.50 2.95 12.25 3.65 ;
    END
END NO5X1
MACRO NO5X2
    CLASS CORE ;
    FOREIGN NO5X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  14.25 2.75 14.75 10.55 ;
        RECT  14.25 7.15 14.95 10.55 ;
        RECT  14.25 2.75 15.15 4.40 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  12.45 5.40 13.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  10.05 4.10 10.95 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  5.25 7.70 5.95 11.00 ;
        RECT  6.75 10.10 7.45 11.00 ;
        RECT  8.25 7.55 8.95 11.00 ;
        RECT  12.90 7.30 13.60 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.70 2.00 3.40 3.60 ;
        RECT  5.40 2.00 6.10 3.60 ;
        RECT  10.05 2.00 10.75 3.40 ;
        RECT  12.90 2.00 13.60 4.40 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.65 4.25 1.15 10.55 ;
        RECT  0.45 8.55 1.15 10.55 ;
        RECT  1.35 2.95 2.05 4.75 ;
        RECT  0.65 7.40 2.60 8.10 ;
        RECT  4.05 2.95 4.75 4.75 ;
        RECT  0.65 4.25 6.50 4.75 ;
        RECT  5.80 4.25 6.50 4.95 ;
        RECT  6.95 3.10 7.45 8.15 ;
        RECT  6.75 7.45 7.45 8.15 ;
        RECT  7.75 2.95 8.45 3.65 ;
        RECT  6.95 3.10 8.45 3.65 ;
        RECT  7.90 5.45 8.60 6.15 ;
        RECT  7.75 2.95 9.50 3.45 ;
        RECT  8.80 2.45 9.50 3.45 ;
        RECT  6.95 3.10 9.50 3.45 ;
        RECT  10.60 5.45 11.10 10.05 ;
        RECT  10.60 7.55 11.30 10.05 ;
        RECT  11.40 2.75 11.90 5.95 ;
        RECT  7.90 5.45 11.90 5.95 ;
        RECT  11.40 2.75 12.10 3.45 ;
    END
END NO5X2
MACRO NO5X3
    CLASS CORE ;
    FOREIGN NO5X3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  13.35 7.15 14.05 10.55 ;
        RECT  14.25 2.45 14.75 7.65 ;
        RECT  13.35 7.15 14.75 7.65 ;
        RECT  13.35 9.85 14.95 10.55 ;
        RECT  14.25 2.45 15.15 4.40 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  12.45 5.25 13.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  10.05 4.10 10.95 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.35 3.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  5.05 7.30 5.75 11.00 ;
        RECT  6.55 10.10 7.25 11.00 ;
        RECT  8.05 7.25 8.75 11.00 ;
        RECT  12.00 7.30 12.70 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.70 2.00 3.40 3.60 ;
        RECT  5.40 2.00 6.10 3.60 ;
        RECT  10.05 2.00 10.75 3.40 ;
        RECT  12.90 2.00 13.60 4.40 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.65 4.25 1.15 10.55 ;
        RECT  0.45 8.55 1.15 10.55 ;
        RECT  1.35 2.95 2.05 4.75 ;
        RECT  0.65 7.40 2.40 8.10 ;
        RECT  4.05 2.95 4.75 4.75 ;
        RECT  5.80 4.05 6.50 4.75 ;
        RECT  0.65 4.25 6.50 4.75 ;
        RECT  6.75 5.20 7.25 7.95 ;
        RECT  6.95 3.10 7.25 7.95 ;
        RECT  6.55 7.25 7.25 7.95 ;
        RECT  6.95 3.10 7.45 5.70 ;
        RECT  6.75 5.20 7.45 5.70 ;
        RECT  7.70 6.10 8.40 6.80 ;
        RECT  7.75 2.95 8.45 3.65 ;
        RECT  6.95 3.10 8.45 3.65 ;
        RECT  7.75 2.95 9.50 3.45 ;
        RECT  8.80 2.45 9.50 3.45 ;
        RECT  6.95 3.10 9.50 3.45 ;
        RECT  10.40 6.10 10.90 9.75 ;
        RECT  10.40 7.25 11.10 9.75 ;
        RECT  11.40 2.75 11.90 6.60 ;
        RECT  7.70 6.10 11.90 6.60 ;
        RECT  11.40 2.75 12.10 3.45 ;
    END
END NO5X3
MACRO NO5X4
    CLASS CORE ;
    FOREIGN NO5X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  14.25 2.75 14.75 10.55 ;
        RECT  14.25 7.15 14.95 10.55 ;
        RECT  14.25 2.75 15.15 4.40 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  12.45 5.40 13.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  10.05 4.10 10.95 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  5.25 7.70 5.95 11.00 ;
        RECT  6.75 10.10 7.45 11.00 ;
        RECT  8.25 7.35 8.95 11.00 ;
        RECT  12.90 7.30 13.60 11.00 ;
        RECT  15.60 7.30 16.30 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.70 2.00 3.40 3.60 ;
        RECT  5.40 2.00 6.10 3.60 ;
        RECT  10.05 2.00 10.75 3.40 ;
        RECT  12.90 2.00 13.60 4.40 ;
        RECT  15.60 2.00 16.30 4.40 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.65 4.25 1.15 10.55 ;
        RECT  0.45 8.55 1.15 10.55 ;
        RECT  1.35 2.95 2.05 4.75 ;
        RECT  0.65 7.40 2.60 8.10 ;
        RECT  4.05 2.95 4.75 4.75 ;
        RECT  0.65 4.25 6.50 4.75 ;
        RECT  5.80 4.25 6.50 4.95 ;
        RECT  6.95 3.10 7.45 8.15 ;
        RECT  6.75 7.45 7.45 8.15 ;
        RECT  7.75 2.95 8.45 3.65 ;
        RECT  6.95 3.10 8.45 3.65 ;
        RECT  7.90 5.45 8.60 6.15 ;
        RECT  7.75 2.95 9.50 3.45 ;
        RECT  8.80 2.45 9.50 3.45 ;
        RECT  6.95 3.10 9.50 3.45 ;
        RECT  10.60 5.45 11.10 10.55 ;
        RECT  10.60 7.35 11.30 10.55 ;
        RECT  11.40 2.75 11.90 5.95 ;
        RECT  7.90 5.45 11.90 5.95 ;
        RECT  11.40 2.75 12.10 3.45 ;
    END
END NO5X4
MACRO NO6I1X1
    CLASS CORE ;
    FOREIGN NO6I1X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  18.45 2.65 18.95 8.80 ;
        RECT  18.25 7.15 18.95 8.80 ;
        RECT  18.20 2.65 19.35 3.70 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        RECT  12.85 5.55 14.10 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  10.05 4.10 11.15 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  14.25 4.10 15.15 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.35 7.05 ;
        RECT  5.45 6.35 6.35 7.05 ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.50 1.15 11.00 ;
        RECT  0.45 10.10 2.50 11.00 ;
        RECT  5.65 7.50 6.35 11.00 ;
        RECT  8.50 7.50 9.00 11.00 ;
        RECT  7.20 10.10 9.00 11.00 ;
        RECT  8.50 7.50 9.20 8.20 ;
        RECT  14.30 7.85 15.00 11.00 ;
        RECT  19.60 7.30 20.30 11.00 ;
        RECT  18.70 10.10 20.30 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 2.00 1.20 3.80 ;
        RECT  3.45 2.00 4.15 3.60 ;
        RECT  6.15 2.00 6.85 3.65 ;
        RECT  11.30 2.00 12.00 3.60 ;
        RECT  14.00 2.00 14.70 3.60 ;
        RECT  16.85 2.00 17.55 3.65 ;
        RECT  19.85 2.00 20.55 4.70 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  11.80 7.50 12.65 7.90 ;
        RECT  2.00 2.95 2.50 9.10 ;
        RECT  1.80 7.50 2.50 9.10 ;
        RECT  2.00 2.95 2.80 3.65 ;
        RECT  3.30 7.55 4.00 10.55 ;
        RECT  3.35 5.45 4.05 6.15 ;
        RECT  2.00 5.65 4.05 6.15 ;
        RECT  4.50 4.15 5.00 8.05 ;
        RECT  4.80 2.95 5.00 8.05 ;
        RECT  3.30 7.55 5.00 8.05 ;
        RECT  4.80 2.95 5.50 4.65 ;
        RECT  4.50 4.15 7.30 4.65 ;
        RECT  6.60 4.15 7.30 4.85 ;
        RECT  7.35 6.55 7.85 8.10 ;
        RECT  7.15 7.40 7.85 8.10 ;
        RECT  8.40 3.15 8.90 7.05 ;
        RECT  7.35 6.55 10.30 7.05 ;
        RECT  9.45 9.25 10.15 10.30 ;
        RECT  9.50 2.95 10.20 3.65 ;
        RECT  8.40 3.15 10.20 3.65 ;
        RECT  9.80 6.55 10.30 8.20 ;
        RECT  9.80 7.50 10.55 8.20 ;
        RECT  9.80 7.65 11.30 8.20 ;
        RECT  10.80 7.65 11.30 9.30 ;
        RECT  10.80 8.60 11.50 9.30 ;
        RECT  10.55 5.45 12.30 6.15 ;
        RECT  11.95 4.35 12.30 9.30 ;
        RECT  11.80 4.35 12.30 7.90 ;
        RECT  11.95 7.50 12.65 9.30 ;
        RECT  12.65 2.95 13.15 4.85 ;
        RECT  11.80 4.35 13.15 4.85 ;
        RECT  12.65 2.95 13.35 3.65 ;
        RECT  13.25 6.85 13.75 10.30 ;
        RECT  9.45 9.80 13.75 10.30 ;
        RECT  15.35 2.95 16.10 3.65 ;
        RECT  15.60 2.95 16.10 7.35 ;
        RECT  13.25 6.85 17.15 7.35 ;
        RECT  16.65 6.85 17.15 10.50 ;
        RECT  16.65 7.50 17.35 10.50 ;
    END
END NO6I1X1
MACRO NO6I1X2
    CLASS CORE ;
    FOREIGN NO6I1X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  18.20 2.65 18.95 4.25 ;
        RECT  18.45 2.65 18.95 10.55 ;
        RECT  18.25 7.15 18.95 10.55 ;
        RECT  18.20 2.65 19.35 3.70 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        RECT  12.85 5.55 14.10 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  10.05 4.10 11.15 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  14.25 4.10 15.15 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.35 7.05 ;
        RECT  5.45 6.35 6.35 7.05 ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.50 1.15 11.00 ;
        RECT  0.45 10.10 2.50 11.00 ;
        RECT  5.65 7.50 6.35 11.00 ;
        RECT  8.50 7.50 9.00 11.00 ;
        RECT  7.20 10.10 9.00 11.00 ;
        RECT  8.50 7.50 9.20 8.20 ;
        RECT  14.30 7.85 15.00 11.00 ;
        RECT  19.60 7.30 20.30 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 2.00 1.20 3.80 ;
        RECT  3.45 2.00 4.15 3.60 ;
        RECT  6.15 2.00 6.85 3.65 ;
        RECT  11.30 2.00 12.00 3.60 ;
        RECT  14.00 2.00 14.70 3.60 ;
        RECT  16.85 2.00 17.55 4.25 ;
        RECT  19.85 2.00 20.55 4.70 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  11.80 7.50 12.65 7.90 ;
        RECT  2.00 2.95 2.50 9.10 ;
        RECT  1.80 7.50 2.50 9.10 ;
        RECT  2.00 2.95 2.80 3.65 ;
        RECT  3.30 7.55 4.00 10.55 ;
        RECT  3.35 5.45 4.05 6.15 ;
        RECT  2.00 5.65 4.05 6.15 ;
        RECT  4.50 4.15 5.00 8.05 ;
        RECT  4.80 2.95 5.00 8.05 ;
        RECT  3.30 7.55 5.00 8.05 ;
        RECT  4.80 2.95 5.50 4.65 ;
        RECT  4.50 4.15 7.30 4.65 ;
        RECT  6.60 4.15 7.30 4.85 ;
        RECT  7.35 6.55 7.85 8.10 ;
        RECT  7.15 7.40 7.85 8.10 ;
        RECT  8.40 3.15 8.90 7.05 ;
        RECT  7.35 6.55 10.30 7.05 ;
        RECT  9.45 9.25 10.15 10.30 ;
        RECT  9.50 2.95 10.20 3.65 ;
        RECT  8.40 3.15 10.20 3.65 ;
        RECT  9.80 6.55 10.30 8.20 ;
        RECT  9.80 7.50 10.55 8.20 ;
        RECT  9.80 7.65 11.30 8.20 ;
        RECT  10.80 7.65 11.30 9.30 ;
        RECT  10.80 8.60 11.50 9.30 ;
        RECT  10.55 5.45 12.30 6.15 ;
        RECT  11.95 4.35 12.30 9.30 ;
        RECT  11.80 4.35 12.30 7.90 ;
        RECT  11.95 7.50 12.65 9.30 ;
        RECT  12.65 2.95 13.15 4.85 ;
        RECT  11.80 4.35 13.15 4.85 ;
        RECT  12.65 2.95 13.35 3.65 ;
        RECT  13.25 6.85 13.75 10.30 ;
        RECT  9.45 9.80 13.75 10.30 ;
        RECT  15.35 2.95 16.10 3.65 ;
        RECT  15.60 2.95 16.10 7.35 ;
        RECT  13.25 6.85 17.15 7.35 ;
        RECT  16.65 6.85 17.15 10.50 ;
        RECT  16.65 7.50 17.35 10.50 ;
    END
END NO6I1X2
MACRO NO6I1X4
    CLASS CORE ;
    FOREIGN NO6I1X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  18.25 2.65 18.95 4.25 ;
        RECT  18.45 2.65 18.95 6.30 ;
        RECT  18.45 5.40 19.35 6.30 ;
        RECT  18.45 5.80 20.10 6.30 ;
        RECT  19.60 5.80 20.10 10.55 ;
        RECT  19.60 7.15 20.30 10.55 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        RECT  12.85 5.55 14.10 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  10.05 4.10 11.15 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  14.25 4.10 15.15 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.35 7.05 ;
        RECT  5.45 6.35 6.35 7.05 ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.50 1.15 11.00 ;
        RECT  0.45 10.10 2.50 11.00 ;
        RECT  5.65 7.50 6.35 11.00 ;
        RECT  8.50 7.50 9.00 11.00 ;
        RECT  7.20 10.10 9.00 11.00 ;
        RECT  8.50 7.50 9.20 8.20 ;
        RECT  14.30 7.85 15.00 11.00 ;
        RECT  18.25 7.30 18.95 11.00 ;
        RECT  20.95 7.30 21.65 11.00 ;
        RECT  0.00 11.00 22.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 2.00 1.20 3.80 ;
        RECT  3.45 2.00 4.15 3.60 ;
        RECT  6.15 2.00 6.85 3.65 ;
        RECT  11.30 2.00 12.00 3.60 ;
        RECT  14.00 2.00 14.70 3.60 ;
        RECT  16.85 2.00 17.55 4.25 ;
        RECT  19.60 2.00 20.30 4.25 ;
        RECT  21.25 2.00 21.95 4.25 ;
        RECT  0.00 0.00 22.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  11.80 7.50 12.65 7.90 ;
        RECT  2.00 2.95 2.50 9.10 ;
        RECT  1.80 7.50 2.50 9.10 ;
        RECT  2.00 2.95 2.80 3.65 ;
        RECT  3.30 7.55 4.00 10.55 ;
        RECT  3.35 5.45 4.05 6.15 ;
        RECT  2.00 5.65 4.05 6.15 ;
        RECT  4.50 4.15 5.00 8.05 ;
        RECT  4.80 2.95 5.00 8.05 ;
        RECT  3.30 7.55 5.00 8.05 ;
        RECT  4.80 2.95 5.50 4.65 ;
        RECT  4.50 4.15 7.30 4.65 ;
        RECT  6.60 4.15 7.30 4.85 ;
        RECT  7.35 6.55 7.85 8.10 ;
        RECT  7.15 7.40 7.85 8.10 ;
        RECT  8.40 3.15 8.90 7.05 ;
        RECT  7.35 6.55 10.30 7.05 ;
        RECT  9.45 9.25 10.15 10.30 ;
        RECT  9.50 2.95 10.20 3.65 ;
        RECT  8.40 3.15 10.20 3.65 ;
        RECT  9.80 6.55 10.30 8.20 ;
        RECT  9.80 7.50 10.55 8.20 ;
        RECT  9.80 7.65 11.30 8.20 ;
        RECT  10.80 7.65 11.30 9.30 ;
        RECT  10.80 8.60 11.50 9.30 ;
        RECT  10.55 5.45 12.30 6.15 ;
        RECT  11.95 4.35 12.30 9.30 ;
        RECT  11.80 4.35 12.30 7.90 ;
        RECT  11.95 7.50 12.65 9.30 ;
        RECT  12.65 2.95 13.15 4.85 ;
        RECT  11.80 4.35 13.15 4.85 ;
        RECT  12.65 2.95 13.35 3.65 ;
        RECT  13.25 6.85 13.75 10.30 ;
        RECT  9.45 9.80 13.75 10.30 ;
        RECT  15.35 2.95 16.10 3.65 ;
        RECT  15.60 2.95 16.10 7.35 ;
        RECT  13.25 6.85 17.15 7.35 ;
        RECT  16.65 6.85 17.15 10.50 ;
        RECT  16.65 7.50 17.35 10.50 ;
    END
END NO6I1X4
MACRO NO6I2X1
    CLASS CORE ;
    FOREIGN NO6I2X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  17.05 2.80 17.95 3.70 ;
        RECT  17.05 3.20 18.70 3.70 ;
        RECT  18.20 3.20 18.70 8.80 ;
        RECT  18.20 7.20 18.90 8.80 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        RECT  11.45 5.55 12.75 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.90 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  12.85 4.10 14.10 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 3.05 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.15 2.50 11.00 ;
        RECT  4.80 7.45 5.35 11.00 ;
        RECT  4.65 9.10 5.35 11.00 ;
        RECT  4.80 7.45 5.50 8.15 ;
        RECT  7.50 7.55 8.00 11.00 ;
        RECT  7.50 7.55 8.20 8.25 ;
        RECT  12.90 7.85 13.60 11.00 ;
        RECT  16.85 7.20 17.55 11.00 ;
        RECT  16.85 10.10 19.15 11.00 ;
        RECT  0.00 11.00 19.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.00 2.00 2.70 4.40 ;
        RECT  2.00 2.00 4.50 2.80 ;
        RECT  5.50 2.00 6.20 2.80 ;
        RECT  10.35 2.00 11.05 3.60 ;
        RECT  13.05 2.00 13.75 3.60 ;
        RECT  15.75 2.00 16.45 3.65 ;
        RECT  0.00 0.00 19.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  10.40 7.50 11.25 8.00 ;
        RECT  0.30 2.45 1.00 3.15 ;
        RECT  0.45 2.45 0.95 9.80 ;
        RECT  0.45 2.45 1.00 4.45 ;
        RECT  0.45 8.15 1.15 9.80 ;
        RECT  0.45 3.75 1.35 4.45 ;
        RECT  1.40 7.00 2.10 7.70 ;
        RECT  1.40 7.20 4.00 7.70 ;
        RECT  3.50 3.95 4.00 9.80 ;
        RECT  3.30 9.10 4.00 9.80 ;
        RECT  4.35 3.75 5.05 4.45 ;
        RECT  3.50 3.95 5.05 4.45 ;
        RECT  6.35 6.60 6.85 8.15 ;
        RECT  6.15 7.45 6.85 8.15 ;
        RECT  6.90 2.90 7.40 7.10 ;
        RECT  6.35 6.60 9.35 7.10 ;
        RECT  8.40 5.45 9.10 6.15 ;
        RECT  8.45 9.80 9.15 10.55 ;
        RECT  8.85 6.60 9.35 8.25 ;
        RECT  8.85 7.55 9.90 8.25 ;
        RECT  8.85 2.70 9.55 3.40 ;
        RECT  6.90 2.90 9.55 3.40 ;
        RECT  9.40 7.55 9.90 9.30 ;
        RECT  9.40 8.60 10.10 9.30 ;
        RECT  8.40 5.65 10.90 6.15 ;
        RECT  10.55 4.35 10.90 9.30 ;
        RECT  10.40 4.35 10.90 8.00 ;
        RECT  10.55 7.50 11.25 9.30 ;
        RECT  11.70 2.95 12.20 4.85 ;
        RECT  10.40 4.35 12.20 4.85 ;
        RECT  11.85 6.85 12.35 10.30 ;
        RECT  8.45 9.80 12.35 10.30 ;
        RECT  11.70 2.95 12.40 3.65 ;
        RECT  14.40 2.95 15.15 3.65 ;
        RECT  14.65 2.95 15.15 7.35 ;
        RECT  11.85 6.85 15.95 7.35 ;
        RECT  15.25 6.85 15.95 10.00 ;
    END
END NO6I2X1
MACRO NO6I2X2
    CLASS CORE ;
    FOREIGN NO6I2X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  17.05 2.65 17.95 3.70 ;
        RECT  17.25 2.65 17.95 4.25 ;
        RECT  17.25 3.75 18.70 4.25 ;
        RECT  18.20 3.75 18.70 10.55 ;
        RECT  18.20 7.15 18.90 10.55 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        RECT  11.45 5.55 12.75 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.90 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  12.85 4.10 14.10 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 3.05 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.15 2.50 11.00 ;
        RECT  4.80 7.45 5.35 11.00 ;
        RECT  4.65 9.10 5.35 11.00 ;
        RECT  4.80 7.45 5.50 8.15 ;
        RECT  7.50 7.55 8.00 11.00 ;
        RECT  7.50 7.55 8.20 8.25 ;
        RECT  12.90 7.85 13.60 11.00 ;
        RECT  16.85 7.30 17.55 11.00 ;
        RECT  0.00 11.00 19.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.00 2.00 2.70 4.40 ;
        RECT  2.00 2.00 4.50 2.80 ;
        RECT  5.50 2.00 6.20 2.80 ;
        RECT  10.35 2.00 11.05 3.60 ;
        RECT  13.05 2.00 13.75 3.60 ;
        RECT  15.90 2.00 16.60 4.25 ;
        RECT  0.00 0.00 19.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  10.40 7.50 11.25 8.00 ;
        RECT  0.30 2.45 1.00 3.15 ;
        RECT  0.45 2.45 0.95 9.80 ;
        RECT  0.45 2.45 1.00 4.45 ;
        RECT  0.45 8.15 1.15 9.80 ;
        RECT  0.45 3.75 1.35 4.45 ;
        RECT  1.40 7.00 2.10 7.70 ;
        RECT  1.40 7.20 4.00 7.70 ;
        RECT  3.50 3.95 4.00 9.80 ;
        RECT  3.30 9.10 4.00 9.80 ;
        RECT  4.35 3.75 5.05 4.45 ;
        RECT  3.50 3.95 5.05 4.45 ;
        RECT  6.35 6.60 6.85 8.15 ;
        RECT  6.15 7.45 6.85 8.15 ;
        RECT  6.90 2.90 7.40 7.10 ;
        RECT  6.35 6.60 9.35 7.10 ;
        RECT  8.40 5.45 9.10 6.15 ;
        RECT  8.45 9.80 9.15 10.55 ;
        RECT  8.85 6.60 9.35 8.25 ;
        RECT  8.85 7.55 9.90 8.25 ;
        RECT  8.85 2.70 9.55 3.40 ;
        RECT  6.90 2.90 9.55 3.40 ;
        RECT  9.40 7.55 9.90 9.30 ;
        RECT  9.40 8.60 10.10 9.30 ;
        RECT  8.40 5.65 10.90 6.15 ;
        RECT  10.55 4.35 10.90 9.30 ;
        RECT  10.40 4.35 10.90 8.00 ;
        RECT  10.55 7.50 11.25 9.30 ;
        RECT  11.70 2.95 12.20 4.85 ;
        RECT  10.40 4.35 12.20 4.85 ;
        RECT  11.85 6.85 12.35 10.30 ;
        RECT  8.45 9.80 12.35 10.30 ;
        RECT  11.70 2.95 12.40 3.65 ;
        RECT  14.40 2.95 15.15 3.65 ;
        RECT  14.65 2.95 15.15 7.35 ;
        RECT  11.85 6.85 15.95 7.35 ;
        RECT  15.25 6.85 15.95 10.00 ;
    END
END NO6I2X2
MACRO NO6I2X4
    CLASS CORE ;
    FOREIGN NO6I2X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  17.25 2.65 17.95 4.25 ;
        RECT  17.45 2.65 17.95 6.30 ;
        RECT  17.05 5.40 17.95 6.30 ;
        RECT  17.05 5.80 18.70 6.30 ;
        RECT  18.20 5.80 18.70 10.55 ;
        RECT  18.20 7.15 18.90 10.55 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        RECT  11.45 5.55 12.75 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.90 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  12.85 4.10 14.10 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 3.05 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.15 2.50 11.00 ;
        RECT  4.80 7.45 5.35 11.00 ;
        RECT  4.65 9.10 5.35 11.00 ;
        RECT  4.80 7.45 5.50 8.15 ;
        RECT  7.50 7.55 8.00 11.00 ;
        RECT  7.50 7.55 8.20 8.25 ;
        RECT  12.90 7.85 13.60 11.00 ;
        RECT  16.85 7.30 17.55 11.00 ;
        RECT  19.55 7.30 20.25 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.00 2.00 2.70 4.40 ;
        RECT  2.00 2.00 4.50 2.80 ;
        RECT  5.50 2.00 6.20 2.80 ;
        RECT  10.35 2.00 11.05 3.60 ;
        RECT  13.05 2.00 13.75 3.60 ;
        RECT  15.90 2.00 16.60 4.25 ;
        RECT  18.60 2.00 19.30 4.25 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  10.40 7.50 11.25 8.00 ;
        RECT  0.30 2.45 1.00 3.15 ;
        RECT  0.45 2.45 0.95 9.80 ;
        RECT  0.45 2.45 1.00 4.45 ;
        RECT  0.45 8.15 1.15 9.80 ;
        RECT  0.45 3.75 1.35 4.45 ;
        RECT  1.40 7.00 2.10 7.70 ;
        RECT  1.40 7.20 4.00 7.70 ;
        RECT  3.50 3.95 4.00 9.80 ;
        RECT  3.30 9.10 4.00 9.80 ;
        RECT  4.35 3.75 5.05 4.45 ;
        RECT  3.50 3.95 5.05 4.45 ;
        RECT  6.35 6.60 6.85 8.15 ;
        RECT  6.15 7.45 6.85 8.15 ;
        RECT  6.90 2.90 7.40 7.10 ;
        RECT  6.35 6.60 9.35 7.10 ;
        RECT  8.40 5.45 9.10 6.15 ;
        RECT  8.45 9.80 9.15 10.55 ;
        RECT  8.85 6.60 9.35 8.25 ;
        RECT  8.85 7.55 9.90 8.25 ;
        RECT  8.85 2.70 9.55 3.40 ;
        RECT  6.90 2.90 9.55 3.40 ;
        RECT  9.40 7.55 9.90 9.30 ;
        RECT  9.40 8.60 10.10 9.30 ;
        RECT  8.40 5.65 10.90 6.15 ;
        RECT  10.55 4.35 10.90 9.30 ;
        RECT  10.40 4.35 10.90 8.00 ;
        RECT  10.55 7.50 11.25 9.30 ;
        RECT  11.70 2.95 12.20 4.85 ;
        RECT  10.40 4.35 12.20 4.85 ;
        RECT  11.85 6.85 12.35 10.30 ;
        RECT  8.45 9.80 12.35 10.30 ;
        RECT  11.70 2.95 12.40 3.65 ;
        RECT  14.40 2.95 15.15 3.65 ;
        RECT  14.65 2.95 15.15 7.35 ;
        RECT  11.85 6.85 15.95 7.35 ;
        RECT  15.25 6.85 15.95 10.00 ;
    END
END NO6I2X4
MACRO NO6I3X1
    CLASS CORE ;
    FOREIGN NO6I3X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  19.85 2.80 20.35 8.80 ;
        RECT  19.85 7.20 20.55 8.80 ;
        RECT  19.85 2.80 20.75 3.70 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        RECT  11.45 5.55 12.75 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.90 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  12.85 4.10 14.05 5.00 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  18.15 5.40 19.35 6.30 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 3.05 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.15 2.50 11.00 ;
        RECT  4.80 7.45 5.35 11.00 ;
        RECT  4.65 9.10 5.35 11.00 ;
        RECT  4.80 7.45 5.50 8.15 ;
        RECT  7.50 7.55 8.00 11.00 ;
        RECT  7.50 7.55 8.20 8.25 ;
        RECT  12.90 7.85 13.60 11.00 ;
        RECT  18.50 7.30 19.20 11.00 ;
        RECT  17.15 10.55 20.55 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.00 2.00 2.70 4.40 ;
        RECT  1.65 2.00 4.15 2.80 ;
        RECT  5.10 2.00 5.80 2.40 ;
        RECT  10.10 2.00 10.80 3.60 ;
        RECT  12.80 2.00 13.50 3.60 ;
        RECT  15.50 2.00 16.20 3.60 ;
        RECT  18.50 2.00 19.20 3.65 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  10.40 7.50 11.25 8.00 ;
        RECT  0.30 2.45 1.00 3.15 ;
        RECT  0.45 2.45 0.95 9.80 ;
        RECT  0.45 2.45 1.00 4.45 ;
        RECT  0.45 8.15 1.15 9.80 ;
        RECT  0.45 3.75 1.35 4.45 ;
        RECT  1.40 7.00 2.10 7.70 ;
        RECT  1.40 7.20 4.00 7.70 ;
        RECT  3.50 4.00 4.00 9.80 ;
        RECT  3.30 9.10 4.00 9.80 ;
        RECT  4.35 3.80 5.05 4.50 ;
        RECT  3.50 4.00 5.05 4.50 ;
        RECT  6.35 6.60 6.85 8.15 ;
        RECT  6.15 7.45 6.85 8.15 ;
        RECT  6.90 2.65 7.40 7.10 ;
        RECT  6.35 6.60 9.35 7.10 ;
        RECT  8.40 5.45 9.10 6.15 ;
        RECT  8.45 9.80 9.15 10.55 ;
        RECT  8.60 2.45 9.30 3.15 ;
        RECT  6.90 2.65 9.30 3.15 ;
        RECT  8.85 6.60 9.35 8.25 ;
        RECT  8.85 7.55 9.90 8.25 ;
        RECT  9.40 7.55 9.90 9.30 ;
        RECT  9.40 8.60 10.10 9.30 ;
        RECT  8.40 5.65 10.90 6.15 ;
        RECT  10.55 4.35 10.90 9.30 ;
        RECT  10.40 4.35 10.90 8.00 ;
        RECT  10.55 7.50 11.25 9.30 ;
        RECT  11.45 2.95 11.95 4.85 ;
        RECT  10.40 4.35 11.95 4.85 ;
        RECT  11.45 2.95 12.15 3.65 ;
        RECT  11.85 6.85 12.35 10.30 ;
        RECT  8.45 9.80 12.35 10.30 ;
        RECT  14.15 2.95 15.00 3.65 ;
        RECT  14.50 2.95 15.00 7.35 ;
        RECT  11.85 6.85 15.95 7.35 ;
        RECT  15.25 6.85 15.95 10.00 ;
        RECT  15.45 5.55 16.15 6.25 ;
        RECT  15.45 5.75 17.65 6.25 ;
        RECT  17.15 2.95 17.65 8.80 ;
        RECT  17.15 2.95 17.85 3.65 ;
        RECT  17.15 7.20 17.85 8.80 ;
    END
END NO6I3X1
MACRO NO6I3X2
    CLASS CORE ;
    FOREIGN NO6I3X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  19.85 2.75 20.35 10.55 ;
        RECT  19.85 2.75 20.55 4.35 ;
        RECT  19.85 7.15 20.55 10.55 ;
        RECT  19.85 2.75 20.75 3.70 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        RECT  11.45 5.55 12.75 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.90 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  12.85 4.10 14.05 5.00 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  18.15 5.40 19.35 6.30 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 3.05 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.15 2.50 11.00 ;
        RECT  4.80 7.45 5.35 11.00 ;
        RECT  4.65 9.10 5.35 11.00 ;
        RECT  4.80 7.45 5.50 8.15 ;
        RECT  7.50 7.55 8.00 11.00 ;
        RECT  7.50 7.55 8.20 8.25 ;
        RECT  12.90 7.85 13.60 11.00 ;
        RECT  16.80 10.20 17.50 11.00 ;
        RECT  18.50 7.30 19.20 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.00 2.00 2.70 4.40 ;
        RECT  1.65 2.00 4.15 2.80 ;
        RECT  5.10 2.00 5.80 2.40 ;
        RECT  10.10 2.00 10.80 3.60 ;
        RECT  12.80 2.00 13.50 3.60 ;
        RECT  15.50 2.00 16.20 3.60 ;
        RECT  18.50 2.00 19.20 4.35 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  10.40 7.50 11.25 8.00 ;
        RECT  0.30 2.45 1.00 3.15 ;
        RECT  0.45 2.45 0.95 9.80 ;
        RECT  0.45 2.45 1.00 4.45 ;
        RECT  0.45 8.15 1.15 9.80 ;
        RECT  0.45 3.75 1.35 4.45 ;
        RECT  1.40 7.00 2.10 7.70 ;
        RECT  1.40 7.20 4.00 7.70 ;
        RECT  3.50 4.00 4.00 9.80 ;
        RECT  3.30 9.10 4.00 9.80 ;
        RECT  4.35 3.80 5.05 4.50 ;
        RECT  3.50 4.00 5.05 4.50 ;
        RECT  6.35 6.60 6.85 8.15 ;
        RECT  6.15 7.45 6.85 8.15 ;
        RECT  6.90 2.65 7.40 7.10 ;
        RECT  6.35 6.60 9.35 7.10 ;
        RECT  8.40 5.45 9.10 6.15 ;
        RECT  8.45 9.80 9.15 10.55 ;
        RECT  8.60 2.45 9.30 3.15 ;
        RECT  6.90 2.65 9.30 3.15 ;
        RECT  8.85 6.60 9.35 8.25 ;
        RECT  8.85 7.55 9.90 8.25 ;
        RECT  9.40 7.55 9.90 9.30 ;
        RECT  9.40 8.60 10.10 9.30 ;
        RECT  8.40 5.65 10.90 6.15 ;
        RECT  10.55 4.35 10.90 9.30 ;
        RECT  10.40 4.35 10.90 8.00 ;
        RECT  10.55 7.50 11.25 9.30 ;
        RECT  11.45 2.95 11.95 4.85 ;
        RECT  10.40 4.35 11.95 4.85 ;
        RECT  11.45 2.95 12.15 3.65 ;
        RECT  11.85 6.85 12.35 10.30 ;
        RECT  8.45 9.80 12.35 10.30 ;
        RECT  14.15 2.95 15.00 3.65 ;
        RECT  14.50 2.95 15.00 7.35 ;
        RECT  11.85 6.85 15.95 7.35 ;
        RECT  15.25 6.85 15.95 10.00 ;
        RECT  15.45 5.55 16.15 6.25 ;
        RECT  15.45 5.75 17.50 6.25 ;
        RECT  17.00 2.95 17.50 8.85 ;
        RECT  17.00 2.95 17.70 3.65 ;
        RECT  17.00 7.15 17.70 8.85 ;
    END
END NO6I3X2
MACRO NO6I3X4
    CLASS CORE ;
    FOREIGN NO6I3X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  19.85 2.75 20.35 10.55 ;
        RECT  19.85 2.75 20.55 4.35 ;
        RECT  19.85 7.15 20.55 10.55 ;
        RECT  19.85 2.75 20.75 3.70 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        RECT  11.45 5.55 12.75 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.90 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  12.85 4.10 14.05 5.00 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  18.15 5.40 19.35 6.30 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 3.05 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.15 2.50 11.00 ;
        RECT  4.80 7.45 5.35 11.00 ;
        RECT  4.65 9.10 5.35 11.00 ;
        RECT  4.80 7.45 5.50 8.15 ;
        RECT  7.50 7.55 8.00 11.00 ;
        RECT  7.50 7.55 8.20 8.25 ;
        RECT  12.90 7.85 13.60 11.00 ;
        RECT  16.80 10.20 17.50 11.00 ;
        RECT  18.50 7.30 19.20 11.00 ;
        RECT  21.20 7.30 21.90 11.00 ;
        RECT  0.00 11.00 22.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.00 2.00 2.70 4.40 ;
        RECT  1.65 2.00 4.15 2.80 ;
        RECT  5.10 2.00 5.80 2.40 ;
        RECT  10.10 2.00 10.80 3.60 ;
        RECT  12.80 2.00 13.50 3.60 ;
        RECT  15.50 2.00 16.20 3.60 ;
        RECT  18.50 2.00 19.20 4.35 ;
        RECT  21.20 2.00 21.90 4.35 ;
        RECT  0.00 0.00 22.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  10.40 7.50 11.25 8.00 ;
        RECT  0.30 2.45 1.00 3.15 ;
        RECT  0.45 2.45 0.95 9.80 ;
        RECT  0.45 2.45 1.00 4.45 ;
        RECT  0.45 8.15 1.15 9.80 ;
        RECT  0.45 3.75 1.35 4.45 ;
        RECT  1.40 7.00 2.10 7.70 ;
        RECT  1.40 7.20 4.00 7.70 ;
        RECT  3.50 4.00 4.00 9.80 ;
        RECT  3.30 9.10 4.00 9.80 ;
        RECT  4.35 3.80 5.05 4.50 ;
        RECT  3.50 4.00 5.05 4.50 ;
        RECT  6.35 6.60 6.85 8.15 ;
        RECT  6.15 7.45 6.85 8.15 ;
        RECT  6.90 2.65 7.40 7.10 ;
        RECT  6.35 6.60 9.35 7.10 ;
        RECT  8.40 5.45 9.10 6.15 ;
        RECT  8.45 9.80 9.15 10.55 ;
        RECT  8.60 2.45 9.30 3.15 ;
        RECT  6.90 2.65 9.30 3.15 ;
        RECT  8.85 6.60 9.35 8.25 ;
        RECT  8.85 7.55 9.90 8.25 ;
        RECT  9.40 7.55 9.90 9.30 ;
        RECT  9.40 8.60 10.10 9.30 ;
        RECT  8.40 5.65 10.90 6.15 ;
        RECT  10.55 4.35 10.90 9.30 ;
        RECT  10.40 4.35 10.90 8.00 ;
        RECT  10.55 7.50 11.25 9.30 ;
        RECT  11.45 2.95 11.95 4.85 ;
        RECT  10.40 4.35 11.95 4.85 ;
        RECT  11.45 2.95 12.15 3.65 ;
        RECT  11.85 6.85 12.35 10.30 ;
        RECT  8.45 9.80 12.35 10.30 ;
        RECT  14.15 2.95 15.00 3.65 ;
        RECT  14.50 2.95 15.00 7.35 ;
        RECT  11.85 6.85 15.95 7.35 ;
        RECT  15.25 6.85 15.95 10.00 ;
        RECT  15.45 5.55 16.15 6.25 ;
        RECT  15.45 5.75 17.50 6.25 ;
        RECT  17.00 2.95 17.50 8.85 ;
        RECT  17.00 2.95 17.70 3.65 ;
        RECT  17.00 7.15 17.70 8.85 ;
    END
END NO6I3X4
MACRO NO6I4X1
    CLASS CORE ;
    FOREIGN NO6I4X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  19.85 3.75 20.35 8.75 ;
        RECT  19.85 7.15 20.55 8.75 ;
        RECT  19.85 3.75 20.75 5.00 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.60 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.90 5.00 ;
        END
    END E
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  12.85 4.10 13.90 5.00 ;
        END
    END DN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  15.30 6.70 16.55 7.60 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 3.05 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.15 2.50 11.00 ;
        RECT  4.80 7.45 5.35 11.00 ;
        RECT  4.65 9.10 5.35 11.00 ;
        RECT  4.80 7.45 5.50 8.15 ;
        RECT  7.50 7.55 8.00 11.00 ;
        RECT  7.50 7.55 8.20 8.25 ;
        RECT  6.80 10.10 9.40 11.00 ;
        RECT  12.80 8.05 13.50 11.00 ;
        RECT  15.50 8.05 16.20 11.00 ;
        RECT  18.50 7.30 19.20 11.00 ;
        RECT  14.65 10.50 20.55 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.00 2.00 2.70 4.40 ;
        RECT  1.65 2.00 4.15 2.80 ;
        RECT  5.10 2.00 5.80 2.40 ;
        RECT  10.10 2.00 10.80 3.60 ;
        RECT  12.80 2.00 13.50 3.60 ;
        RECT  18.50 2.00 19.20 4.40 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  17.15 3.75 17.85 4.45 ;
        RECT  8.85 7.55 9.80 8.25 ;
        RECT  0.30 2.45 1.00 3.15 ;
        RECT  0.45 2.45 0.95 9.80 ;
        RECT  0.45 2.45 1.00 4.45 ;
        RECT  0.45 8.15 1.15 9.80 ;
        RECT  0.45 3.75 1.35 4.45 ;
        RECT  1.40 7.00 2.10 7.70 ;
        RECT  1.40 7.20 4.00 7.70 ;
        RECT  3.50 4.00 4.00 9.80 ;
        RECT  3.30 9.10 4.00 9.80 ;
        RECT  4.35 3.80 5.05 4.50 ;
        RECT  3.50 4.00 5.05 4.50 ;
        RECT  6.35 6.60 6.85 8.15 ;
        RECT  6.15 7.45 6.85 8.15 ;
        RECT  6.90 2.65 7.40 7.10 ;
        RECT  6.35 6.60 9.35 7.10 ;
        RECT  8.40 5.45 9.10 6.15 ;
        RECT  8.60 2.45 9.30 3.15 ;
        RECT  6.90 2.65 9.30 3.15 ;
        RECT  9.30 6.60 9.35 9.65 ;
        RECT  8.85 6.60 9.35 8.25 ;
        RECT  9.30 7.55 9.80 9.65 ;
        RECT  9.30 8.95 10.00 9.65 ;
        RECT  8.40 5.65 10.95 6.15 ;
        RECT  10.45 4.35 10.95 10.50 ;
        RECT  10.45 7.50 11.15 10.50 ;
        RECT  11.45 2.95 11.95 4.85 ;
        RECT  10.45 4.35 11.95 4.85 ;
        RECT  11.45 2.95 12.15 3.65 ;
        RECT  14.35 5.10 14.85 8.75 ;
        RECT  14.15 8.05 14.85 8.75 ;
        RECT  15.15 2.95 15.85 3.65 ;
        RECT  15.35 2.95 15.85 5.60 ;
        RECT  14.35 5.10 16.90 5.60 ;
        RECT  16.20 5.10 16.90 5.80 ;
        RECT  16.55 2.45 17.65 3.15 ;
        RECT  17.35 2.45 17.65 8.85 ;
        RECT  17.15 2.45 17.65 4.45 ;
        RECT  17.35 3.75 17.85 8.85 ;
        RECT  17.15 7.15 17.85 8.85 ;
    END
END NO6I4X1
MACRO NO6I4X2
    CLASS CORE ;
    FOREIGN NO6I4X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  19.85 2.75 20.35 10.55 ;
        RECT  19.85 2.75 20.55 4.35 ;
        RECT  19.85 7.15 20.55 10.55 ;
        RECT  19.85 2.75 20.75 3.70 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.60 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.90 5.00 ;
        END
    END E
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  12.85 4.10 13.90 5.00 ;
        END
    END DN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  15.30 6.70 16.55 7.60 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 3.05 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.15 2.50 11.00 ;
        RECT  4.80 7.45 5.35 11.00 ;
        RECT  4.65 9.10 5.35 11.00 ;
        RECT  4.80 7.45 5.50 8.15 ;
        RECT  7.50 7.55 8.00 11.00 ;
        RECT  7.50 7.55 8.20 8.25 ;
        RECT  6.80 10.10 9.40 11.00 ;
        RECT  12.80 8.05 13.50 11.00 ;
        RECT  15.50 8.05 16.20 11.00 ;
        RECT  14.65 10.20 17.45 11.00 ;
        RECT  18.50 7.30 19.20 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.00 2.00 2.70 4.40 ;
        RECT  1.65 2.00 4.15 2.80 ;
        RECT  5.10 2.00 5.80 2.40 ;
        RECT  10.10 2.00 10.80 3.60 ;
        RECT  12.80 2.00 13.50 3.60 ;
        RECT  18.50 2.00 19.20 4.35 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  8.85 7.55 9.80 8.25 ;
        RECT  0.30 2.45 1.00 3.15 ;
        RECT  0.45 2.45 0.95 9.80 ;
        RECT  0.45 2.45 1.00 4.45 ;
        RECT  0.45 8.15 1.15 9.80 ;
        RECT  0.45 3.75 1.35 4.45 ;
        RECT  1.40 7.00 2.10 7.70 ;
        RECT  1.40 7.20 4.00 7.70 ;
        RECT  3.50 4.00 4.00 9.80 ;
        RECT  3.30 9.10 4.00 9.80 ;
        RECT  4.35 3.80 5.05 4.50 ;
        RECT  3.50 4.00 5.05 4.50 ;
        RECT  6.35 6.60 6.85 8.15 ;
        RECT  6.15 7.45 6.85 8.15 ;
        RECT  6.90 2.65 7.40 7.10 ;
        RECT  6.35 6.60 9.35 7.10 ;
        RECT  8.40 5.45 9.10 6.15 ;
        RECT  8.60 2.45 9.30 3.15 ;
        RECT  6.90 2.65 9.30 3.15 ;
        RECT  9.30 6.60 9.35 9.65 ;
        RECT  8.85 6.60 9.35 8.25 ;
        RECT  9.30 7.55 9.80 9.65 ;
        RECT  9.30 8.95 10.00 9.65 ;
        RECT  8.40 5.65 10.95 6.15 ;
        RECT  10.45 4.35 10.95 10.50 ;
        RECT  10.45 7.50 11.15 10.50 ;
        RECT  11.45 2.95 11.95 4.85 ;
        RECT  10.45 4.35 11.95 4.85 ;
        RECT  11.45 2.95 12.15 3.65 ;
        RECT  14.35 5.10 14.85 8.75 ;
        RECT  14.15 8.05 14.85 8.75 ;
        RECT  15.15 2.95 15.85 3.65 ;
        RECT  15.35 2.95 15.85 5.60 ;
        RECT  14.35 5.10 16.75 5.60 ;
        RECT  16.05 5.10 16.75 5.80 ;
        RECT  16.65 2.45 17.70 3.15 ;
        RECT  17.00 3.75 17.70 4.45 ;
        RECT  17.20 2.45 17.70 8.85 ;
        RECT  17.00 7.15 17.70 8.85 ;
    END
END NO6I4X2
MACRO NO6I4X4
    CLASS CORE ;
    FOREIGN NO6I4X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  19.85 2.75 20.35 10.55 ;
        RECT  19.85 2.75 20.55 4.45 ;
        RECT  19.85 7.15 20.55 10.55 ;
        RECT  19.85 2.75 20.75 3.70 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.60 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.90 5.00 ;
        END
    END E
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  12.85 4.10 13.90 5.00 ;
        END
    END DN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  15.30 6.70 16.55 7.60 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 3.05 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.15 2.50 11.00 ;
        RECT  4.80 7.45 5.35 11.00 ;
        RECT  4.65 9.10 5.35 11.00 ;
        RECT  4.80 7.45 5.50 8.15 ;
        RECT  7.50 7.55 8.00 11.00 ;
        RECT  7.50 7.55 8.20 8.25 ;
        RECT  6.80 10.10 9.40 11.00 ;
        RECT  12.80 8.05 13.50 11.00 ;
        RECT  15.50 8.05 16.20 11.00 ;
        RECT  14.65 10.20 17.45 11.00 ;
        RECT  18.50 7.30 19.20 11.00 ;
        RECT  21.20 7.30 21.90 11.00 ;
        RECT  0.00 11.00 22.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.00 2.00 2.70 4.40 ;
        RECT  1.65 2.00 4.15 2.80 ;
        RECT  5.10 2.00 5.80 2.40 ;
        RECT  10.10 2.00 10.80 3.60 ;
        RECT  12.80 2.00 13.50 3.60 ;
        RECT  18.50 2.00 19.20 4.45 ;
        RECT  21.20 2.00 21.90 4.45 ;
        RECT  0.00 0.00 22.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  8.85 7.55 9.80 8.25 ;
        RECT  0.30 2.45 1.00 3.15 ;
        RECT  0.45 2.45 0.95 9.80 ;
        RECT  0.45 2.45 1.00 4.45 ;
        RECT  0.45 8.15 1.15 9.80 ;
        RECT  0.45 3.75 1.35 4.45 ;
        RECT  1.40 7.00 2.10 7.70 ;
        RECT  1.40 7.20 4.00 7.70 ;
        RECT  3.50 4.00 4.00 9.80 ;
        RECT  3.30 9.10 4.00 9.80 ;
        RECT  4.35 3.80 5.05 4.50 ;
        RECT  3.50 4.00 5.05 4.50 ;
        RECT  6.35 6.60 6.85 8.15 ;
        RECT  6.15 7.45 6.85 8.15 ;
        RECT  6.90 2.65 7.40 7.10 ;
        RECT  6.35 6.60 9.35 7.10 ;
        RECT  8.40 5.45 9.10 6.15 ;
        RECT  8.60 2.45 9.30 3.15 ;
        RECT  6.90 2.65 9.30 3.15 ;
        RECT  9.30 6.60 9.35 9.65 ;
        RECT  8.85 6.60 9.35 8.25 ;
        RECT  9.30 7.55 9.80 9.65 ;
        RECT  9.30 8.95 10.00 9.65 ;
        RECT  8.40 5.65 10.95 6.15 ;
        RECT  10.45 4.35 10.95 10.50 ;
        RECT  10.45 7.50 11.15 10.50 ;
        RECT  11.45 2.95 11.95 4.85 ;
        RECT  10.45 4.35 11.95 4.85 ;
        RECT  11.45 2.95 12.15 3.65 ;
        RECT  14.35 5.10 14.85 8.75 ;
        RECT  14.15 8.05 14.85 8.75 ;
        RECT  15.15 2.95 15.85 3.65 ;
        RECT  15.35 2.95 15.85 5.60 ;
        RECT  14.35 5.10 16.75 5.60 ;
        RECT  16.05 5.10 16.75 5.80 ;
        RECT  16.65 2.45 17.70 3.15 ;
        RECT  17.00 3.75 17.70 4.45 ;
        RECT  17.20 2.45 17.70 8.85 ;
        RECT  17.00 7.15 17.70 8.85 ;
    END
END NO6I4X4
MACRO NO6I5X1
    CLASS CORE ;
    FOREIGN NO6I5X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  22.65 2.80 23.15 8.75 ;
        RECT  22.65 2.80 23.35 4.40 ;
        RECT  22.65 7.15 23.35 8.75 ;
        RECT  22.65 2.80 23.55 3.70 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.40 6.30 ;
        END
    END F
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.90 6.30 ;
        END
    END EN
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  15.65 4.10 16.70 5.00 ;
        END
    END DN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  18.25 6.70 19.35 7.60 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 3.05 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.15 2.50 11.00 ;
        RECT  4.80 7.45 5.35 11.00 ;
        RECT  4.65 9.10 5.35 11.00 ;
        RECT  4.80 7.45 5.50 8.15 ;
        RECT  7.50 7.55 8.00 11.00 ;
        RECT  7.50 7.55 8.20 8.25 ;
        RECT  6.80 10.10 9.40 11.00 ;
        RECT  12.75 7.60 13.45 11.00 ;
        RECT  15.75 8.15 16.45 11.00 ;
        RECT  18.45 8.15 19.15 11.00 ;
        RECT  21.30 7.30 22.00 11.00 ;
        RECT  0.00 11.00 23.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.00 2.00 2.70 4.40 ;
        RECT  1.60 2.00 4.10 2.65 ;
        RECT  4.90 2.00 5.60 2.40 ;
        RECT  10.10 2.00 10.80 3.05 ;
        RECT  12.80 2.00 13.50 3.05 ;
        RECT  15.75 2.00 16.45 3.60 ;
        RECT  21.30 2.00 22.00 4.40 ;
        RECT  0.00 0.00 23.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  19.95 3.75 20.65 4.45 ;
        RECT  8.85 7.55 9.75 8.25 ;
        RECT  0.30 2.45 1.00 3.15 ;
        RECT  0.45 2.45 0.95 9.80 ;
        RECT  0.45 2.45 1.00 4.45 ;
        RECT  0.45 8.15 1.15 9.80 ;
        RECT  0.45 3.75 1.35 4.45 ;
        RECT  1.40 7.00 2.10 7.70 ;
        RECT  1.40 7.20 4.00 7.70 ;
        RECT  3.50 4.00 4.00 9.80 ;
        RECT  3.30 9.10 4.00 9.80 ;
        RECT  4.35 3.80 5.05 4.50 ;
        RECT  3.50 4.00 5.05 4.50 ;
        RECT  6.35 6.60 6.85 8.15 ;
        RECT  6.15 7.45 6.85 8.15 ;
        RECT  7.00 2.65 7.50 7.10 ;
        RECT  7.95 5.45 8.65 6.15 ;
        RECT  6.35 6.60 9.35 7.10 ;
        RECT  8.40 2.45 9.10 3.15 ;
        RECT  7.00 2.65 9.10 3.15 ;
        RECT  9.25 6.60 9.35 9.65 ;
        RECT  8.85 6.60 9.35 8.25 ;
        RECT  9.25 7.55 9.75 9.65 ;
        RECT  9.40 3.50 9.90 6.15 ;
        RECT  9.25 8.95 9.95 9.65 ;
        RECT  7.95 5.65 10.90 6.15 ;
        RECT  10.40 5.65 10.90 10.50 ;
        RECT  10.35 4.45 11.05 5.15 ;
        RECT  10.40 7.50 11.10 10.50 ;
        RECT  11.45 2.45 11.95 4.00 ;
        RECT  9.40 3.50 11.95 4.00 ;
        RECT  11.45 2.45 12.15 3.15 ;
        RECT  14.15 2.45 14.95 3.15 ;
        RECT  10.35 4.45 14.95 4.95 ;
        RECT  14.45 2.45 14.95 9.20 ;
        RECT  14.25 7.60 14.95 9.20 ;
        RECT  17.30 5.10 17.80 8.85 ;
        RECT  17.10 8.15 17.80 8.85 ;
        RECT  18.10 2.95 18.80 3.65 ;
        RECT  18.30 2.95 18.80 5.60 ;
        RECT  17.30 5.10 19.55 5.60 ;
        RECT  18.85 5.10 19.55 5.80 ;
        RECT  19.45 2.45 20.45 3.15 ;
        RECT  20.15 2.45 20.45 8.85 ;
        RECT  19.95 2.45 20.45 4.45 ;
        RECT  20.15 3.75 20.65 8.85 ;
        RECT  19.95 7.15 20.65 8.85 ;
    END
END NO6I5X1
MACRO NO6I5X2
    CLASS CORE ;
    FOREIGN NO6I5X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  22.65 2.75 23.15 10.55 ;
        RECT  22.65 2.75 23.35 4.35 ;
        RECT  22.65 7.15 23.35 10.55 ;
        RECT  22.65 2.75 23.55 3.70 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.40 6.30 ;
        END
    END F
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.90 6.30 ;
        END
    END EN
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  15.65 4.10 16.70 5.00 ;
        END
    END DN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  18.10 6.70 19.35 7.60 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 3.05 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.15 2.50 11.00 ;
        RECT  4.80 7.45 5.35 11.00 ;
        RECT  4.65 9.10 5.35 11.00 ;
        RECT  4.80 7.45 5.50 8.15 ;
        RECT  7.50 7.55 8.00 11.00 ;
        RECT  7.50 7.55 8.20 8.25 ;
        RECT  6.80 10.10 9.40 11.00 ;
        RECT  12.75 7.60 13.45 11.00 ;
        RECT  15.60 8.15 16.30 11.00 ;
        RECT  18.30 8.15 19.00 11.00 ;
        RECT  14.50 10.20 19.70 11.00 ;
        RECT  21.30 7.30 22.00 11.00 ;
        RECT  0.00 11.00 23.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.00 2.00 2.70 4.40 ;
        RECT  1.60 2.00 4.10 2.65 ;
        RECT  4.90 2.00 5.60 2.40 ;
        RECT  10.10 2.00 10.80 3.05 ;
        RECT  12.80 2.00 13.50 3.05 ;
        RECT  15.65 2.00 16.35 3.60 ;
        RECT  21.30 2.00 22.00 4.35 ;
        RECT  0.00 0.00 23.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  19.80 3.75 20.50 4.45 ;
        RECT  8.85 7.55 9.75 8.25 ;
        RECT  0.30 2.45 1.00 3.15 ;
        RECT  0.45 2.45 0.95 9.80 ;
        RECT  0.45 2.45 1.00 4.45 ;
        RECT  0.45 8.15 1.15 9.80 ;
        RECT  0.45 3.75 1.35 4.45 ;
        RECT  1.40 7.00 2.10 7.70 ;
        RECT  1.40 7.20 4.00 7.70 ;
        RECT  3.50 4.00 4.00 9.80 ;
        RECT  3.30 9.10 4.00 9.80 ;
        RECT  4.35 3.80 5.05 4.50 ;
        RECT  3.50 4.00 5.05 4.50 ;
        RECT  6.35 6.60 6.85 8.15 ;
        RECT  6.15 7.45 6.85 8.15 ;
        RECT  7.00 2.65 7.50 7.10 ;
        RECT  7.95 5.45 8.65 6.15 ;
        RECT  6.35 6.60 9.35 7.10 ;
        RECT  8.40 2.45 9.10 3.15 ;
        RECT  7.00 2.65 9.10 3.15 ;
        RECT  9.25 6.60 9.35 9.65 ;
        RECT  8.85 6.60 9.35 8.25 ;
        RECT  9.25 7.55 9.75 9.65 ;
        RECT  9.40 3.50 9.90 6.15 ;
        RECT  9.25 8.95 9.95 9.65 ;
        RECT  7.95 5.65 10.90 6.15 ;
        RECT  10.40 5.65 10.90 10.50 ;
        RECT  10.35 4.45 11.05 5.15 ;
        RECT  10.40 7.50 11.10 10.50 ;
        RECT  11.45 2.45 11.95 4.00 ;
        RECT  9.40 3.50 11.95 4.00 ;
        RECT  11.45 2.45 12.15 3.15 ;
        RECT  14.15 2.45 14.85 3.15 ;
        RECT  10.35 4.45 14.85 4.95 ;
        RECT  14.35 2.45 14.85 9.20 ;
        RECT  14.10 7.60 14.85 9.20 ;
        RECT  17.15 5.10 17.65 8.85 ;
        RECT  16.95 8.15 17.65 8.85 ;
        RECT  18.00 2.95 18.70 3.65 ;
        RECT  18.20 2.95 18.70 5.60 ;
        RECT  17.15 5.10 19.55 5.60 ;
        RECT  18.85 5.10 19.55 5.80 ;
        RECT  19.45 2.45 20.30 3.15 ;
        RECT  20.00 2.45 20.30 8.85 ;
        RECT  19.80 2.45 20.30 4.45 ;
        RECT  20.00 3.75 20.50 8.85 ;
        RECT  19.80 7.15 20.50 8.85 ;
    END
END NO6I5X2
MACRO NO6I5X4
    CLASS CORE ;
    FOREIGN NO6I5X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 25.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  22.65 2.75 23.15 10.55 ;
        RECT  22.65 2.75 23.35 4.35 ;
        RECT  22.65 7.15 23.35 10.55 ;
        RECT  22.65 2.75 23.55 3.70 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.40 6.30 ;
        END
    END F
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.90 6.30 ;
        END
    END EN
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  15.65 4.10 16.70 5.00 ;
        END
    END DN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  18.10 6.70 19.35 7.60 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 3.05 6.30 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.15 2.50 11.00 ;
        RECT  4.80 7.45 5.35 11.00 ;
        RECT  4.65 9.10 5.35 11.00 ;
        RECT  4.80 7.45 5.50 8.15 ;
        RECT  7.50 7.55 8.00 11.00 ;
        RECT  7.50 7.55 8.20 8.25 ;
        RECT  6.80 10.10 9.40 11.00 ;
        RECT  12.75 7.60 13.45 11.00 ;
        RECT  15.60 8.15 16.30 11.00 ;
        RECT  18.30 8.15 19.00 11.00 ;
        RECT  14.50 10.20 19.70 11.00 ;
        RECT  21.30 7.30 22.00 11.00 ;
        RECT  24.00 7.30 24.70 11.00 ;
        RECT  0.00 11.00 25.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.00 2.00 2.70 4.40 ;
        RECT  1.60 2.00 4.10 2.65 ;
        RECT  4.90 2.00 5.60 2.40 ;
        RECT  10.10 2.00 10.80 3.05 ;
        RECT  12.80 2.00 13.50 3.05 ;
        RECT  15.65 2.00 16.35 3.60 ;
        RECT  21.30 2.00 22.00 4.35 ;
        RECT  24.00 2.00 24.70 4.35 ;
        RECT  0.00 0.00 25.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  19.80 3.75 20.50 4.45 ;
        RECT  8.85 7.55 9.75 8.25 ;
        RECT  0.30 2.45 1.00 3.15 ;
        RECT  0.45 2.45 0.95 9.80 ;
        RECT  0.45 2.45 1.00 4.45 ;
        RECT  0.45 8.15 1.15 9.80 ;
        RECT  0.45 3.75 1.35 4.45 ;
        RECT  1.40 7.00 2.10 7.70 ;
        RECT  1.40 7.20 4.00 7.70 ;
        RECT  3.50 4.00 4.00 9.80 ;
        RECT  3.30 9.10 4.00 9.80 ;
        RECT  4.35 3.80 5.05 4.50 ;
        RECT  3.50 4.00 5.05 4.50 ;
        RECT  6.35 6.60 6.85 8.15 ;
        RECT  6.15 7.45 6.85 8.15 ;
        RECT  7.00 2.65 7.50 7.10 ;
        RECT  7.95 5.45 8.65 6.15 ;
        RECT  6.35 6.60 9.35 7.10 ;
        RECT  8.40 2.45 9.10 3.15 ;
        RECT  7.00 2.65 9.10 3.15 ;
        RECT  9.25 6.60 9.35 9.65 ;
        RECT  8.85 6.60 9.35 8.25 ;
        RECT  9.25 7.55 9.75 9.65 ;
        RECT  9.40 3.50 9.90 6.15 ;
        RECT  9.25 8.95 9.95 9.65 ;
        RECT  7.95 5.65 10.90 6.15 ;
        RECT  10.40 5.65 10.90 10.50 ;
        RECT  10.35 4.45 11.05 5.15 ;
        RECT  10.40 7.50 11.10 10.50 ;
        RECT  11.45 2.45 11.95 4.00 ;
        RECT  9.40 3.50 11.95 4.00 ;
        RECT  11.45 2.45 12.15 3.15 ;
        RECT  14.15 2.45 14.85 3.15 ;
        RECT  10.35 4.45 14.85 4.95 ;
        RECT  14.35 2.45 14.85 9.20 ;
        RECT  14.10 7.60 14.85 9.20 ;
        RECT  17.15 5.10 17.65 8.85 ;
        RECT  16.95 8.15 17.65 8.85 ;
        RECT  18.00 2.95 18.70 3.65 ;
        RECT  18.20 2.95 18.70 5.60 ;
        RECT  17.15 5.10 19.55 5.60 ;
        RECT  18.85 5.10 19.55 5.80 ;
        RECT  19.45 2.45 20.30 3.15 ;
        RECT  20.00 2.45 20.30 8.85 ;
        RECT  19.80 2.45 20.30 4.45 ;
        RECT  20.00 3.75 20.50 8.85 ;
        RECT  19.80 7.15 20.50 8.85 ;
    END
END NO6I5X4
MACRO NO6X1
    CLASS CORE ;
    FOREIGN NO6X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  15.40 3.00 16.10 3.70 ;
        RECT  15.60 3.00 16.10 7.20 ;
        RECT  15.60 6.70 17.30 7.20 ;
        RECT  16.80 6.70 17.30 9.30 ;
        RECT  16.80 7.70 17.50 9.30 ;
        RECT  16.80 8.00 17.95 8.90 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.30 ;
        RECT  10.05 5.55 11.30 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  7.25 4.10 8.35 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  11.45 4.10 12.50 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.55 7.05 ;
        RECT  2.25 6.35 3.55 7.05 ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.95 9.25 3.65 11.00 ;
        RECT  4.25 8.65 4.75 11.00 ;
        RECT  5.30 7.60 5.80 9.15 ;
        RECT  4.25 8.65 5.80 9.15 ;
        RECT  5.30 7.60 6.00 8.30 ;
        RECT  11.50 7.85 12.20 11.00 ;
        RECT  15.45 7.70 16.15 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.30 ;
        RECT  3.15 2.00 3.85 3.35 ;
        RECT  8.65 2.00 9.35 3.60 ;
        RECT  11.35 2.00 12.05 3.60 ;
        RECT  14.05 2.00 14.75 3.65 ;
        RECT  17.05 2.00 17.75 4.65 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  9.00 7.50 9.85 7.90 ;
        RECT  0.45 7.55 1.15 10.05 ;
        RECT  1.25 5.45 1.75 8.05 ;
        RECT  1.60 2.65 1.75 8.05 ;
        RECT  0.45 7.55 1.75 8.05 ;
        RECT  1.60 2.65 1.95 5.95 ;
        RECT  1.25 5.45 1.95 5.95 ;
        RECT  1.60 2.65 2.10 5.90 ;
        RECT  1.25 5.45 2.10 5.90 ;
        RECT  1.60 2.65 2.50 3.35 ;
        RECT  1.60 3.85 4.20 4.35 ;
        RECT  3.50 3.85 4.20 4.55 ;
        RECT  4.35 6.65 4.85 8.20 ;
        RECT  3.95 7.50 4.85 8.20 ;
        RECT  5.20 9.60 5.90 10.30 ;
        RECT  5.50 2.90 6.00 7.15 ;
        RECT  4.35 6.65 7.15 7.15 ;
        RECT  6.65 6.65 7.15 8.30 ;
        RECT  6.50 2.70 7.20 3.40 ;
        RECT  5.50 2.90 7.20 3.40 ;
        RECT  6.65 7.60 7.35 8.30 ;
        RECT  6.65 7.75 8.50 8.30 ;
        RECT  7.65 5.60 8.35 6.30 ;
        RECT  8.00 7.75 8.50 9.30 ;
        RECT  8.00 8.60 8.70 9.30 ;
        RECT  7.65 5.80 9.50 6.30 ;
        RECT  9.15 4.35 9.50 9.30 ;
        RECT  9.00 4.35 9.50 7.90 ;
        RECT  9.15 7.50 9.85 9.30 ;
        RECT  10.00 2.95 10.50 4.85 ;
        RECT  9.00 4.35 10.50 4.85 ;
        RECT  10.00 2.95 10.70 3.65 ;
        RECT  10.45 6.85 10.95 10.30 ;
        RECT  5.20 9.80 10.95 10.30 ;
        RECT  12.70 2.95 13.45 3.65 ;
        RECT  12.95 2.95 13.45 7.35 ;
        RECT  10.45 6.85 14.35 7.35 ;
        RECT  13.85 6.85 14.35 10.00 ;
        RECT  13.85 7.50 14.55 10.00 ;
    END
END NO6X1
MACRO NO6X2
    CLASS CORE ;
    FOREIGN NO6X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  15.40 2.65 16.15 4.25 ;
        RECT  15.65 2.65 16.15 10.55 ;
        RECT  15.45 7.15 16.15 10.55 ;
        RECT  15.40 2.65 16.55 3.70 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.30 ;
        RECT  10.05 5.55 11.30 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  7.25 4.10 8.35 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  11.45 4.10 12.35 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.55 7.05 ;
        RECT  2.25 6.35 3.55 7.05 ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 7.50 3.50 11.00 ;
        RECT  5.50 7.50 6.00 11.00 ;
        RECT  5.50 7.50 6.20 8.20 ;
        RECT  11.50 7.85 12.20 11.00 ;
        RECT  16.80 7.30 17.50 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.30 ;
        RECT  3.15 2.00 3.85 3.35 ;
        RECT  8.50 2.00 9.20 3.60 ;
        RECT  11.20 2.00 11.90 3.60 ;
        RECT  14.05 2.00 14.75 4.25 ;
        RECT  17.05 2.00 17.75 4.70 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  9.00 7.50 9.85 7.90 ;
        RECT  0.45 7.55 1.15 10.05 ;
        RECT  1.25 5.45 1.75 8.05 ;
        RECT  1.60 2.65 1.75 8.05 ;
        RECT  0.45 7.55 1.75 8.05 ;
        RECT  1.60 2.65 1.95 5.95 ;
        RECT  1.25 5.45 1.95 5.95 ;
        RECT  1.60 2.65 2.10 5.90 ;
        RECT  1.25 5.45 2.10 5.90 ;
        RECT  1.60 2.65 2.50 3.35 ;
        RECT  1.60 3.85 4.30 4.35 ;
        RECT  3.60 3.85 4.30 4.55 ;
        RECT  4.35 6.55 4.85 8.10 ;
        RECT  4.15 7.40 4.85 8.10 ;
        RECT  5.50 2.90 6.00 7.05 ;
        RECT  4.35 6.55 7.35 7.05 ;
        RECT  6.45 9.25 7.15 10.30 ;
        RECT  6.50 2.70 7.20 3.40 ;
        RECT  5.50 2.90 7.20 3.40 ;
        RECT  6.85 6.55 7.35 8.20 ;
        RECT  6.85 7.50 7.55 8.20 ;
        RECT  6.85 7.65 8.50 8.20 ;
        RECT  8.00 7.65 8.50 9.30 ;
        RECT  8.00 8.60 8.70 9.30 ;
        RECT  7.75 5.60 9.50 6.30 ;
        RECT  9.15 4.35 9.50 9.30 ;
        RECT  9.00 4.35 9.50 7.90 ;
        RECT  9.15 7.50 9.85 9.30 ;
        RECT  9.85 2.95 10.35 4.85 ;
        RECT  9.00 4.35 10.35 4.85 ;
        RECT  9.85 2.95 10.55 3.65 ;
        RECT  10.45 6.85 10.95 10.30 ;
        RECT  6.45 9.80 10.95 10.30 ;
        RECT  12.55 2.95 13.30 3.65 ;
        RECT  12.80 2.95 13.30 7.35 ;
        RECT  10.45 6.85 14.35 7.35 ;
        RECT  13.85 6.85 14.35 10.00 ;
        RECT  13.85 7.50 14.55 10.00 ;
    END
END NO6X2
MACRO NO6X3
    CLASS CORE ;
    FOREIGN NO6X3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  15.40 2.65 16.15 4.25 ;
        RECT  15.45 7.15 16.15 10.55 ;
        RECT  15.65 2.65 16.15 10.55 ;
        RECT  14.55 9.85 16.15 10.55 ;
        RECT  15.40 2.65 16.55 3.70 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  7.25 4.10 8.35 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  11.45 4.10 12.35 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.55 7.15 ;
        RECT  2.25 6.45 3.55 7.15 ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 7.60 3.50 11.00 ;
        RECT  5.35 7.60 5.85 11.00 ;
        RECT  5.35 7.60 6.20 8.30 ;
        RECT  11.05 7.75 11.75 11.00 ;
        RECT  16.80 7.20 17.50 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.30 ;
        RECT  3.15 2.00 3.85 3.35 ;
        RECT  8.50 2.00 9.20 3.60 ;
        RECT  11.20 2.00 11.90 3.60 ;
        RECT  14.05 2.00 14.75 4.25 ;
        RECT  17.05 2.00 17.75 4.70 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 7.65 1.15 10.15 ;
        RECT  1.25 5.45 1.75 8.15 ;
        RECT  0.45 7.65 1.75 8.15 ;
        RECT  1.80 2.65 2.30 5.95 ;
        RECT  1.25 5.45 2.30 5.95 ;
        RECT  1.80 2.65 2.50 4.35 ;
        RECT  1.80 3.85 4.30 4.35 ;
        RECT  3.60 3.85 4.30 4.55 ;
        RECT  4.35 6.55 4.85 8.20 ;
        RECT  4.15 7.50 4.85 8.20 ;
        RECT  5.50 2.90 6.00 7.05 ;
        RECT  4.35 6.55 7.35 7.05 ;
        RECT  6.30 9.35 7.00 10.30 ;
        RECT  6.50 2.70 7.20 3.40 ;
        RECT  5.50 2.90 7.20 3.40 ;
        RECT  6.85 6.55 7.35 8.30 ;
        RECT  6.85 7.60 8.05 8.30 ;
        RECT  7.55 7.60 8.05 9.35 ;
        RECT  7.55 8.65 8.25 9.35 ;
        RECT  7.75 5.60 9.40 6.30 ;
        RECT  8.90 4.35 9.40 9.20 ;
        RECT  8.70 7.40 9.40 9.20 ;
        RECT  9.85 2.95 10.35 4.85 ;
        RECT  8.90 4.35 10.35 4.85 ;
        RECT  10.00 6.75 10.50 10.30 ;
        RECT  6.30 9.80 10.50 10.30 ;
        RECT  9.85 2.95 10.55 3.65 ;
        RECT  12.55 2.95 13.30 3.65 ;
        RECT  12.80 2.95 13.30 7.25 ;
        RECT  10.00 6.75 13.90 7.25 ;
        RECT  13.40 6.75 13.90 9.00 ;
        RECT  13.40 7.40 14.10 9.00 ;
    END
END NO6X3
MACRO NO6X4
    CLASS CORE ;
    FOREIGN NO6X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  15.40 2.65 16.10 4.25 ;
        RECT  15.60 2.65 16.10 5.90 ;
        RECT  15.60 5.40 17.95 5.90 ;
        RECT  16.80 5.40 17.50 10.55 ;
        RECT  16.80 5.40 17.95 6.30 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.30 ;
        RECT  10.05 5.55 11.30 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  7.25 4.10 8.35 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  11.45 4.10 12.35 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.55 7.05 ;
        RECT  2.25 6.35 3.55 7.05 ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 7.50 3.50 11.00 ;
        RECT  5.50 7.50 6.00 11.00 ;
        RECT  5.50 7.50 6.20 8.20 ;
        RECT  11.50 7.85 12.20 11.00 ;
        RECT  15.45 7.30 16.15 11.00 ;
        RECT  18.15 7.30 18.85 11.00 ;
        RECT  0.00 11.00 19.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.30 ;
        RECT  3.15 2.00 3.85 3.35 ;
        RECT  8.50 2.00 9.20 3.60 ;
        RECT  11.20 2.00 11.90 3.60 ;
        RECT  14.05 2.00 14.75 4.25 ;
        RECT  16.75 2.00 17.45 4.25 ;
        RECT  18.40 2.00 19.10 4.70 ;
        RECT  0.00 0.00 19.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  9.00 7.50 9.85 7.90 ;
        RECT  0.45 7.55 1.15 10.05 ;
        RECT  1.25 5.45 1.75 8.05 ;
        RECT  1.60 2.65 1.75 8.05 ;
        RECT  0.45 7.55 1.75 8.05 ;
        RECT  1.60 2.65 1.95 5.95 ;
        RECT  1.25 5.45 1.95 5.95 ;
        RECT  1.60 2.65 2.10 5.90 ;
        RECT  1.25 5.45 2.10 5.90 ;
        RECT  1.60 2.65 2.50 3.35 ;
        RECT  1.60 3.85 4.30 4.35 ;
        RECT  3.60 3.85 4.30 4.55 ;
        RECT  4.35 6.55 4.85 8.10 ;
        RECT  4.15 7.40 4.85 8.10 ;
        RECT  5.50 2.90 6.00 7.05 ;
        RECT  4.35 6.55 7.35 7.05 ;
        RECT  6.45 9.25 7.15 10.30 ;
        RECT  6.50 2.70 7.20 3.40 ;
        RECT  5.50 2.90 7.20 3.40 ;
        RECT  6.85 6.55 7.35 8.20 ;
        RECT  6.85 7.50 8.50 8.20 ;
        RECT  8.00 7.50 8.50 9.30 ;
        RECT  8.00 8.60 8.70 9.30 ;
        RECT  7.75 5.60 9.50 6.30 ;
        RECT  9.15 4.35 9.50 9.30 ;
        RECT  9.00 4.35 9.50 7.90 ;
        RECT  9.15 7.50 9.85 9.30 ;
        RECT  9.85 2.95 10.35 4.85 ;
        RECT  9.00 4.35 10.35 4.85 ;
        RECT  9.85 2.95 10.55 3.65 ;
        RECT  10.45 6.85 10.95 10.30 ;
        RECT  6.45 9.80 10.95 10.30 ;
        RECT  12.55 2.95 13.30 3.65 ;
        RECT  12.80 2.95 13.30 7.35 ;
        RECT  10.45 6.85 14.55 7.35 ;
        RECT  13.85 6.85 14.55 10.00 ;
    END
END NO6X4
MACRO NO7X1
    CLASS CORE ;
    FOREIGN NO7X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.25 3.95 0.75 10.20 ;
        RECT  1.10 2.55 1.60 4.45 ;
        RECT  0.25 3.95 1.60 4.45 ;
        RECT  1.10 2.55 1.80 3.25 ;
        RECT  0.25 9.25 1.85 10.20 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  15.60 5.35 16.55 6.15 ;
        RECT  14.90 5.45 16.55 6.15 ;
        RECT  15.65 5.35 16.55 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.40 19.35 6.35 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  13.80 4.50 14.30 5.55 ;
        RECT  13.80 4.50 15.15 5.00 ;
        RECT  14.25 4.10 14.30 5.55 ;
        RECT  13.60 4.85 14.30 5.55 ;
        RECT  14.25 4.10 15.15 5.00 ;
        RECT  13.60 4.85 15.15 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  12.15 4.80 12.35 6.30 ;
        RECT  11.45 5.40 12.35 6.30 ;
        RECT  12.15 4.80 12.85 5.90 ;
        RECT  11.45 5.40 12.85 5.90 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.05 9.85 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.15 10.75 1.85 11.00 ;
        RECT  1.20 7.95 1.90 8.65 ;
        RECT  1.20 8.15 2.85 8.65 ;
        RECT  2.35 8.15 2.85 11.00 ;
        RECT  5.75 7.40 6.45 11.00 ;
        RECT  8.60 7.50 9.30 8.20 ;
        RECT  8.80 7.50 9.30 9.05 ;
        RECT  8.80 8.55 10.05 9.05 ;
        RECT  9.55 8.55 10.05 11.00 ;
        RECT  13.85 6.50 14.55 11.00 ;
        RECT  18.45 9.55 19.15 11.00 ;
        RECT  0.00 11.00 19.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.45 2.00 3.15 3.25 ;
        RECT  5.15 2.00 5.85 3.25 ;
        RECT  11.35 2.00 12.05 3.40 ;
        RECT  14.05 2.00 14.75 3.45 ;
        RECT  16.75 2.00 17.45 3.45 ;
        RECT  0.00 0.00 19.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  7.90 6.90 11.20 6.95 ;
        RECT  6.95 7.45 7.95 7.95 ;
        RECT  3.75 2.55 3.85 10.45 ;
        RECT  3.35 4.10 3.85 10.45 ;
        RECT  3.35 7.45 4.10 10.45 ;
        RECT  3.75 2.55 4.25 4.60 ;
        RECT  3.75 2.55 4.50 3.25 ;
        RECT  3.35 4.10 6.20 4.60 ;
        RECT  5.50 4.10 6.20 4.80 ;
        RECT  7.25 2.75 7.45 10.20 ;
        RECT  6.95 2.75 7.45 7.95 ;
        RECT  7.25 7.45 7.75 10.20 ;
        RECT  6.95 9.30 7.75 10.20 ;
        RECT  7.25 7.45 7.95 8.15 ;
        RECT  6.95 9.70 9.05 10.20 ;
        RECT  7.90 6.25 8.60 6.95 ;
        RECT  8.35 9.70 9.05 10.40 ;
        RECT  8.50 2.55 9.20 3.25 ;
        RECT  6.95 2.75 9.20 3.25 ;
        RECT  10.00 2.75 10.85 3.45 ;
        RECT  10.35 2.75 10.85 7.60 ;
        RECT  10.35 6.90 11.20 7.60 ;
        RECT  10.50 2.75 10.85 10.30 ;
        RECT  7.90 6.45 10.85 6.95 ;
        RECT  10.50 6.90 11.20 10.30 ;
        RECT  12.70 2.75 13.20 4.35 ;
        RECT  10.35 3.85 13.20 4.35 ;
        RECT  12.70 2.75 13.40 3.45 ;
        RECT  15.40 2.75 16.10 3.45 ;
        RECT  15.60 2.75 16.10 4.40 ;
        RECT  17.00 3.90 17.15 10.35 ;
        RECT  16.40 7.25 17.15 10.35 ;
        RECT  17.00 3.90 17.50 7.80 ;
        RECT  16.40 7.25 17.50 7.80 ;
        RECT  15.60 3.90 18.65 4.40 ;
        RECT  17.95 3.90 18.65 4.60 ;
    END
END NO7X1
MACRO NO7X2
    CLASS CORE ;
    FOREIGN NO7X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.70 4.10 1.20 10.50 ;
        RECT  0.95 2.75 1.20 10.50 ;
        RECT  0.50 7.10 1.20 10.50 ;
        RECT  0.95 2.75 1.65 5.00 ;
        RECT  0.25 4.10 1.65 5.00 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  14.90 5.45 16.55 6.15 ;
        RECT  15.60 5.35 16.55 6.35 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.40 19.35 6.35 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  13.80 4.10 15.15 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  11.45 4.10 12.40 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  8.65 3.90 9.85 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.85 7.15 2.55 11.00 ;
        RECT  5.75 7.70 6.45 11.00 ;
        RECT  8.60 7.50 10.05 8.20 ;
        RECT  9.55 7.50 10.05 11.00 ;
        RECT  13.85 6.50 14.55 11.00 ;
        RECT  18.45 9.55 19.15 11.00 ;
        RECT  0.00 11.00 19.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.30 2.00 3.00 4.35 ;
        RECT  5.15 2.00 5.85 3.45 ;
        RECT  11.40 2.00 12.10 3.40 ;
        RECT  14.15 2.00 14.85 3.45 ;
        RECT  16.85 2.00 17.55 3.45 ;
        RECT  0.00 0.00 19.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.80 2.75 4.50 3.45 ;
        RECT  3.40 6.75 4.10 10.45 ;
        RECT  4.00 2.75 4.50 4.60 ;
        RECT  4.00 4.10 6.30 4.60 ;
        RECT  5.50 4.10 6.30 4.80 ;
        RECT  5.80 4.10 6.30 7.25 ;
        RECT  3.40 6.75 6.30 7.25 ;
        RECT  6.95 2.75 7.45 10.20 ;
        RECT  6.95 9.30 7.65 10.20 ;
        RECT  6.95 7.45 7.95 8.15 ;
        RECT  6.95 9.70 9.05 10.20 ;
        RECT  8.15 6.00 8.85 6.70 ;
        RECT  8.35 9.70 9.05 10.40 ;
        RECT  8.50 2.55 9.20 3.25 ;
        RECT  6.95 2.75 9.20 3.25 ;
        RECT  10.00 2.75 10.80 3.45 ;
        RECT  10.50 2.75 10.80 10.30 ;
        RECT  10.30 2.75 10.80 6.70 ;
        RECT  10.50 6.20 11.20 10.30 ;
        RECT  12.85 2.75 13.35 6.70 ;
        RECT  8.15 6.20 13.35 6.70 ;
        RECT  12.80 2.75 13.50 3.45 ;
        RECT  15.50 2.75 16.20 3.45 ;
        RECT  15.70 2.75 16.20 4.40 ;
        RECT  17.00 3.90 17.15 10.55 ;
        RECT  16.40 7.55 17.15 10.55 ;
        RECT  17.00 3.90 17.50 8.10 ;
        RECT  16.40 7.55 17.50 8.10 ;
        RECT  18.00 2.45 18.50 4.40 ;
        RECT  15.70 3.90 18.50 4.40 ;
        RECT  18.00 2.45 18.70 3.15 ;
    END
END NO7X2
MACRO NO7X3
    CLASS CORE ;
    FOREIGN NO7X3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  2.10 4.10 2.60 9.75 ;
        RECT  2.50 3.05 2.60 9.75 ;
        RECT  1.90 7.25 2.60 9.75 ;
        RECT  2.50 3.05 3.00 5.00 ;
        RECT  1.65 4.10 3.00 5.00 ;
        RECT  2.50 3.05 3.20 3.75 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  16.30 5.45 17.95 6.15 ;
        RECT  17.00 5.35 17.95 6.35 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.40 20.75 6.35 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  15.20 4.10 16.55 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  12.85 4.10 13.80 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  10.05 3.90 11.25 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.55 7.25 1.25 11.00 ;
        RECT  3.25 7.25 3.95 11.00 ;
        RECT  7.15 7.70 7.85 11.00 ;
        RECT  10.00 7.50 11.45 8.20 ;
        RECT  10.95 7.50 11.45 11.00 ;
        RECT  15.25 6.50 15.95 11.00 ;
        RECT  19.85 9.55 20.55 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.15 2.00 1.85 3.45 ;
        RECT  3.85 2.00 4.55 3.45 ;
        RECT  6.55 2.00 7.25 3.45 ;
        RECT  12.80 2.00 13.50 3.40 ;
        RECT  15.55 2.00 16.25 3.45 ;
        RECT  18.25 2.00 18.95 3.45 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  5.20 2.75 5.90 3.45 ;
        RECT  4.80 6.75 5.50 10.45 ;
        RECT  5.40 2.75 5.90 4.60 ;
        RECT  5.40 4.10 7.70 4.60 ;
        RECT  6.90 4.10 7.70 4.80 ;
        RECT  7.20 4.10 7.70 7.25 ;
        RECT  4.80 6.75 7.70 7.25 ;
        RECT  8.35 2.75 8.85 10.20 ;
        RECT  8.35 9.30 9.05 10.20 ;
        RECT  8.35 7.45 9.35 8.15 ;
        RECT  8.35 9.70 10.45 10.20 ;
        RECT  9.55 6.00 10.25 6.70 ;
        RECT  9.75 9.70 10.45 10.40 ;
        RECT  9.90 2.55 10.60 3.25 ;
        RECT  8.35 2.75 10.60 3.25 ;
        RECT  11.40 2.75 12.20 3.45 ;
        RECT  11.90 2.75 12.20 10.30 ;
        RECT  11.70 2.75 12.20 6.70 ;
        RECT  11.90 6.20 12.60 10.30 ;
        RECT  14.25 2.75 14.75 6.70 ;
        RECT  9.55 6.20 14.75 6.70 ;
        RECT  14.20 2.75 14.90 3.45 ;
        RECT  16.90 2.75 17.60 3.45 ;
        RECT  17.10 2.75 17.60 4.40 ;
        RECT  18.40 3.90 18.55 10.55 ;
        RECT  17.80 7.55 18.55 10.55 ;
        RECT  18.40 3.90 18.90 8.10 ;
        RECT  17.80 7.55 18.90 8.10 ;
        RECT  19.40 2.45 19.90 4.40 ;
        RECT  17.10 3.90 19.90 4.40 ;
        RECT  19.40 2.45 20.10 3.15 ;
    END
END NO7X3
MACRO NO7X4
    CLASS CORE ;
    FOREIGN NO7X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  2.35 2.80 2.60 10.55 ;
        RECT  1.90 5.40 2.60 10.55 ;
        RECT  2.35 2.80 2.85 6.30 ;
        RECT  1.65 5.40 2.85 6.30 ;
        RECT  2.35 2.80 3.05 4.40 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  16.30 5.45 17.95 6.15 ;
        RECT  17.00 5.35 17.95 6.35 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.40 20.75 6.35 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  15.20 4.10 16.55 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  12.85 4.10 13.80 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  10.05 3.90 11.25 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.55 7.25 1.25 11.00 ;
        RECT  3.25 7.25 3.95 11.00 ;
        RECT  7.15 7.70 7.85 11.00 ;
        RECT  10.00 7.50 11.45 8.20 ;
        RECT  10.95 7.50 11.45 11.00 ;
        RECT  15.25 6.50 15.95 11.00 ;
        RECT  19.85 9.55 20.55 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.00 2.00 1.70 4.40 ;
        RECT  3.70 2.00 4.40 4.40 ;
        RECT  6.55 2.00 7.25 3.45 ;
        RECT  12.80 2.00 13.50 3.40 ;
        RECT  15.55 2.00 16.25 3.45 ;
        RECT  18.25 2.00 18.95 3.45 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  5.20 2.75 5.90 3.45 ;
        RECT  4.80 6.75 5.50 10.45 ;
        RECT  5.40 2.75 5.90 4.60 ;
        RECT  5.40 4.10 7.70 4.60 ;
        RECT  6.90 4.10 7.70 4.80 ;
        RECT  7.20 4.10 7.70 7.25 ;
        RECT  4.80 6.75 7.70 7.25 ;
        RECT  8.35 2.75 8.85 10.20 ;
        RECT  8.35 9.30 9.05 10.20 ;
        RECT  8.35 7.45 9.35 8.15 ;
        RECT  8.35 9.70 10.45 10.20 ;
        RECT  9.55 6.00 10.25 6.70 ;
        RECT  9.75 9.70 10.45 10.40 ;
        RECT  9.90 2.55 10.60 3.25 ;
        RECT  8.35 2.75 10.60 3.25 ;
        RECT  11.40 2.75 12.20 3.45 ;
        RECT  11.90 2.75 12.20 10.30 ;
        RECT  11.70 2.75 12.20 6.70 ;
        RECT  11.90 6.20 12.60 10.30 ;
        RECT  14.25 2.75 14.75 6.70 ;
        RECT  9.55 6.20 14.75 6.70 ;
        RECT  14.20 2.75 14.90 3.45 ;
        RECT  16.90 2.75 17.60 3.45 ;
        RECT  17.10 2.75 17.60 4.40 ;
        RECT  18.40 3.90 18.55 10.55 ;
        RECT  17.80 7.55 18.55 10.55 ;
        RECT  18.40 3.90 18.90 8.10 ;
        RECT  17.80 7.55 18.90 8.10 ;
        RECT  19.40 2.45 19.90 4.40 ;
        RECT  17.10 3.90 19.90 4.40 ;
        RECT  19.40 2.45 20.10 3.15 ;
    END
END NO7X4
MACRO NO8X1
    CLASS CORE ;
    FOREIGN NO8X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  9.75 3.25 10.25 9.35 ;
        RECT  9.55 7.70 10.25 9.35 ;
        RECT  9.60 3.25 10.30 3.95 ;
        RECT  9.75 5.40 10.95 6.30 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  3.00 5.25 3.95 6.30 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  4.10 4.00 4.90 4.70 ;
        RECT  4.40 4.00 4.90 6.30 ;
        RECT  4.40 5.40 5.35 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  5.80 4.50 6.50 6.30 ;
        RECT  5.80 5.40 6.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.30 8.15 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.25 17.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.40 19.35 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.60 7.10 4.30 11.00 ;
        RECT  10.90 7.05 11.60 11.00 ;
        RECT  10.90 7.05 13.30 7.75 ;
        RECT  15.45 7.20 16.15 11.00 ;
        RECT  15.45 10.45 17.20 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 3.40 ;
        RECT  3.65 2.00 4.35 3.45 ;
        RECT  6.50 2.00 7.20 3.10 ;
        RECT  10.95 2.00 11.65 3.90 ;
        RECT  15.80 2.00 16.50 3.05 ;
        RECT  18.50 2.00 19.20 3.10 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.40 4.00 2.10 4.70 ;
        RECT  1.60 4.00 2.10 10.05 ;
        RECT  1.25 7.15 2.10 10.05 ;
        RECT  2.30 2.75 2.80 4.50 ;
        RECT  0.40 4.00 2.80 4.50 ;
        RECT  2.30 2.75 3.00 3.45 ;
        RECT  5.00 2.75 5.85 3.45 ;
        RECT  5.35 2.75 5.85 4.05 ;
        RECT  6.95 7.00 7.65 10.55 ;
        RECT  5.35 3.55 9.10 4.05 ;
        RECT  8.60 2.75 8.70 7.50 ;
        RECT  8.00 2.75 8.70 4.05 ;
        RECT  8.60 3.55 9.10 7.50 ;
        RECT  6.95 7.00 9.10 7.50 ;
        RECT  6.95 9.85 9.10 10.55 ;
        RECT  12.45 2.45 12.95 5.10 ;
        RECT  11.30 4.40 12.95 5.10 ;
        RECT  12.40 8.65 13.10 9.35 ;
        RECT  12.45 2.45 13.15 3.15 ;
        RECT  11.30 4.60 14.45 5.10 ;
        RECT  13.95 4.60 14.45 9.15 ;
        RECT  12.40 8.65 14.45 9.15 ;
        RECT  13.95 7.05 14.65 7.80 ;
        RECT  14.95 4.20 15.65 4.95 ;
        RECT  17.15 2.45 17.85 3.15 ;
        RECT  17.35 2.45 17.85 4.70 ;
        RECT  14.95 4.20 20.35 4.70 ;
        RECT  18.80 7.10 20.55 7.80 ;
        RECT  19.85 2.45 20.35 10.45 ;
        RECT  19.85 2.45 20.55 3.15 ;
        RECT  19.85 7.10 20.55 10.45 ;
    END
END NO8X1
MACRO NO8X2
    CLASS CORE ;
    FOREIGN NO8X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  9.75 2.45 10.25 10.55 ;
        RECT  9.55 7.10 10.25 10.55 ;
        RECT  9.60 2.45 10.30 4.05 ;
        RECT  9.75 5.40 10.95 6.30 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  3.00 5.25 3.95 6.30 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  4.10 4.00 4.90 4.70 ;
        RECT  4.40 4.00 4.90 6.30 ;
        RECT  4.40 5.40 5.35 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  5.80 4.50 6.50 6.30 ;
        RECT  5.80 5.40 6.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.30 8.15 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.25 17.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.40 19.35 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.60 7.10 4.30 11.00 ;
        RECT  10.90 7.15 11.60 11.00 ;
        RECT  10.90 7.15 13.30 7.85 ;
        RECT  15.45 7.20 16.15 11.00 ;
        RECT  15.45 10.45 17.20 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 3.40 ;
        RECT  3.65 2.00 4.35 3.45 ;
        RECT  6.50 2.00 7.20 3.10 ;
        RECT  10.95 2.00 11.65 3.90 ;
        RECT  15.80 2.00 16.50 3.05 ;
        RECT  18.50 2.00 19.20 3.10 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.40 4.00 2.10 4.70 ;
        RECT  1.60 4.00 2.10 10.05 ;
        RECT  1.25 7.15 2.10 10.05 ;
        RECT  2.30 2.75 2.80 4.50 ;
        RECT  0.40 4.00 2.80 4.50 ;
        RECT  2.30 2.75 3.00 3.45 ;
        RECT  5.00 2.75 5.85 3.45 ;
        RECT  5.35 2.75 5.85 4.05 ;
        RECT  6.95 7.00 7.65 10.55 ;
        RECT  5.35 3.55 9.10 4.05 ;
        RECT  8.60 2.75 8.70 7.50 ;
        RECT  8.00 2.75 8.70 4.05 ;
        RECT  8.60 3.55 9.10 7.50 ;
        RECT  6.95 7.00 9.10 7.50 ;
        RECT  6.95 9.85 9.10 10.55 ;
        RECT  12.45 2.45 12.95 5.10 ;
        RECT  11.30 4.40 12.95 5.10 ;
        RECT  12.40 8.75 13.10 9.45 ;
        RECT  12.45 2.45 13.15 3.15 ;
        RECT  11.30 4.60 14.45 5.10 ;
        RECT  13.95 4.60 14.45 9.25 ;
        RECT  12.40 8.75 14.45 9.25 ;
        RECT  13.95 7.15 14.65 7.90 ;
        RECT  14.95 4.20 15.65 4.95 ;
        RECT  17.15 2.45 17.85 3.15 ;
        RECT  17.35 2.45 17.85 4.70 ;
        RECT  14.95 4.20 20.35 4.70 ;
        RECT  18.80 7.10 20.55 7.80 ;
        RECT  19.85 2.45 20.35 10.45 ;
        RECT  19.85 2.45 20.55 3.15 ;
        RECT  19.85 7.10 20.55 10.45 ;
    END
END NO8X2
MACRO NO8X3
    CLASS CORE ;
    FOREIGN NO8X3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  9.60 2.45 10.30 4.05 ;
        RECT  9.60 7.10 10.30 10.10 ;
        RECT  9.80 2.45 10.30 10.10 ;
        RECT  8.30 9.40 10.30 10.10 ;
        RECT  9.80 5.40 10.95 6.30 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  2.70 5.25 3.95 6.30 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  4.10 4.00 4.90 4.70 ;
        RECT  4.40 4.00 4.90 6.30 ;
        RECT  4.40 5.40 5.35 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  5.80 4.50 6.50 6.30 ;
        RECT  5.80 5.40 6.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.30 8.15 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.25 17.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.40 19.35 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.30 7.10 4.00 11.00 ;
        RECT  10.95 7.10 11.65 11.00 ;
        RECT  9.50 10.75 11.65 11.00 ;
        RECT  12.60 6.95 12.75 7.80 ;
        RECT  10.95 7.10 12.75 7.80 ;
        RECT  12.60 6.95 13.30 7.65 ;
        RECT  10.95 7.10 13.30 7.65 ;
        RECT  15.45 7.20 16.15 11.00 ;
        RECT  15.45 10.45 17.20 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 3.40 ;
        RECT  3.65 2.00 4.35 3.45 ;
        RECT  6.50 2.00 7.20 3.10 ;
        RECT  10.95 2.00 11.65 4.20 ;
        RECT  15.80 2.00 16.50 3.05 ;
        RECT  18.50 2.00 19.20 3.10 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.40 4.00 2.10 4.70 ;
        RECT  1.60 4.00 1.65 10.05 ;
        RECT  0.95 7.15 1.65 10.05 ;
        RECT  1.60 4.00 2.10 7.65 ;
        RECT  0.95 7.15 2.10 7.65 ;
        RECT  2.30 2.75 2.80 4.50 ;
        RECT  0.40 4.00 2.80 4.50 ;
        RECT  2.30 2.75 3.00 3.45 ;
        RECT  5.00 2.75 5.85 3.45 ;
        RECT  5.35 2.75 5.85 4.05 ;
        RECT  6.65 6.75 7.35 9.50 ;
        RECT  5.35 3.55 9.10 4.05 ;
        RECT  6.65 8.20 8.40 8.90 ;
        RECT  8.60 2.75 8.70 7.25 ;
        RECT  8.00 2.75 8.70 4.05 ;
        RECT  8.60 3.55 9.10 7.25 ;
        RECT  6.65 6.75 9.10 7.25 ;
        RECT  12.45 2.45 12.95 5.50 ;
        RECT  11.40 4.80 12.95 5.50 ;
        RECT  12.45 2.45 13.15 3.15 ;
        RECT  12.45 8.60 13.15 9.30 ;
        RECT  11.40 5.00 14.45 5.50 ;
        RECT  13.95 5.00 14.45 9.10 ;
        RECT  12.45 8.60 14.45 9.10 ;
        RECT  13.95 7.00 14.65 7.75 ;
        RECT  14.95 4.20 15.65 4.95 ;
        RECT  17.15 2.45 17.85 3.15 ;
        RECT  17.35 2.45 17.85 4.70 ;
        RECT  14.95 4.20 20.35 4.70 ;
        RECT  18.80 7.10 20.55 7.80 ;
        RECT  19.85 2.45 20.35 10.45 ;
        RECT  19.85 2.45 20.55 3.15 ;
        RECT  19.85 7.10 20.55 10.45 ;
    END
END NO8X3
MACRO NO8X4
    CLASS CORE ;
    FOREIGN NO8X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.95 2.45 11.65 4.05 ;
        RECT  11.15 2.45 11.65 10.55 ;
        RECT  10.95 7.10 11.65 10.55 ;
        RECT  11.15 5.40 12.35 6.30 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  3.00 5.25 3.95 6.30 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  4.10 4.00 4.90 4.70 ;
        RECT  4.40 4.00 4.90 6.30 ;
        RECT  4.40 5.40 5.35 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  5.80 4.50 6.50 6.30 ;
        RECT  5.80 5.40 6.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.30 8.15 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.25 19.35 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.60 7.10 4.30 11.00 ;
        RECT  9.60 7.15 10.30 11.00 ;
        RECT  12.30 7.15 13.00 11.00 ;
        RECT  12.30 7.15 14.70 7.85 ;
        RECT  16.85 7.20 17.55 11.00 ;
        RECT  16.85 10.45 18.60 11.00 ;
        RECT  0.00 11.00 22.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 3.40 ;
        RECT  3.65 2.00 4.35 3.45 ;
        RECT  6.50 2.00 7.20 3.10 ;
        RECT  9.60 2.00 10.30 3.90 ;
        RECT  12.30 2.00 13.00 3.90 ;
        RECT  17.20 2.00 17.90 3.05 ;
        RECT  19.90 2.00 20.60 3.10 ;
        RECT  0.00 0.00 22.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.40 4.00 2.10 4.70 ;
        RECT  1.60 4.00 2.10 10.05 ;
        RECT  1.25 7.15 2.10 10.05 ;
        RECT  2.30 2.75 2.80 4.50 ;
        RECT  0.40 4.00 2.80 4.50 ;
        RECT  2.30 2.75 3.00 3.45 ;
        RECT  5.00 2.75 5.85 3.45 ;
        RECT  5.35 2.75 5.85 4.05 ;
        RECT  6.95 7.00 7.65 10.55 ;
        RECT  5.35 3.55 9.10 4.05 ;
        RECT  8.60 2.75 8.70 7.50 ;
        RECT  8.00 2.75 8.70 4.05 ;
        RECT  8.60 3.55 9.10 7.50 ;
        RECT  6.95 7.00 9.10 7.50 ;
        RECT  6.95 9.85 9.10 10.55 ;
        RECT  13.85 2.45 14.35 5.10 ;
        RECT  12.70 4.40 14.35 5.10 ;
        RECT  13.80 8.75 14.50 9.45 ;
        RECT  13.85 2.45 14.55 3.15 ;
        RECT  12.70 4.60 15.85 5.10 ;
        RECT  15.35 4.60 15.85 9.25 ;
        RECT  13.80 8.75 15.85 9.25 ;
        RECT  15.35 7.15 16.05 7.90 ;
        RECT  16.35 4.20 17.05 4.95 ;
        RECT  18.55 2.45 19.25 3.15 ;
        RECT  18.75 2.45 19.25 4.70 ;
        RECT  16.35 4.20 21.75 4.70 ;
        RECT  20.20 7.10 21.95 7.80 ;
        RECT  21.25 2.45 21.75 10.45 ;
        RECT  21.25 2.45 21.95 3.15 ;
        RECT  21.25 7.10 21.95 10.45 ;
    END
END NO8X4
MACRO OA211X1
    CLASS CORE ;
    FOREIGN OA211X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  7.25 3.05 8.15 3.75 ;
        RECT  7.25 5.40 8.15 6.30 ;
        RECT  7.65 3.05 7.90 10.55 ;
        RECT  7.20 8.75 7.90 10.55 ;
        RECT  7.65 3.05 8.15 9.30 ;
        RECT  7.20 8.75 8.15 9.30 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.55 7.60 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  0.25 6.70 1.15 7.60 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 9.05 3.50 11.00 ;
        RECT  5.85 8.90 6.55 11.00 ;
        RECT  0.00 11.00 8.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  5.70 2.00 6.40 3.75 ;
        RECT  0.00 0.00 8.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 2.55 1.15 4.00 ;
        RECT  0.45 8.10 1.15 10.55 ;
        RECT  1.80 3.55 2.50 4.25 ;
        RECT  2.00 3.55 2.50 5.75 ;
        RECT  2.00 5.25 3.55 5.75 ;
        RECT  0.45 2.55 3.85 3.05 ;
        RECT  3.05 5.25 3.55 8.60 ;
        RECT  3.15 2.55 3.85 4.00 ;
        RECT  0.45 8.10 5.00 8.60 ;
        RECT  4.50 7.75 5.00 10.55 ;
        RECT  4.30 9.85 5.00 10.55 ;
        RECT  4.50 7.75 7.20 8.25 ;
        RECT  6.50 7.55 7.20 8.25 ;
        RECT  0.45 8.10 7.20 8.25 ;
    END
END OA211X1
MACRO OA211X2
    CLASS CORE ;
    FOREIGN OA211X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        RECT  7.00 2.50 7.75 4.20 ;
        RECT  7.65 2.50 7.75 10.55 ;
        RECT  7.25 2.50 7.75 6.30 ;
        RECT  7.65 5.40 7.90 10.55 ;
        RECT  7.20 7.95 7.90 10.55 ;
        RECT  7.65 5.40 8.15 8.70 ;
        RECT  7.20 7.95 8.15 8.70 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.55 7.60 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  0.25 6.70 1.15 7.60 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 9.05 3.50 11.00 ;
        RECT  5.80 7.95 6.55 11.00 ;
        RECT  0.00 11.00 8.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  5.65 2.00 6.35 4.20 ;
        RECT  0.00 0.00 8.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 2.55 1.15 4.00 ;
        RECT  0.45 8.10 1.15 10.55 ;
        RECT  1.80 3.55 2.50 4.25 ;
        RECT  2.00 3.55 2.50 5.75 ;
        RECT  2.00 5.25 3.55 5.75 ;
        RECT  0.45 2.55 3.85 3.05 ;
        RECT  3.05 5.25 3.55 8.60 ;
        RECT  3.15 2.55 3.85 4.00 ;
        RECT  0.45 8.10 5.00 8.60 ;
        RECT  4.50 7.00 5.00 10.55 ;
        RECT  4.30 9.85 5.00 10.55 ;
        RECT  6.50 6.80 7.20 7.50 ;
        RECT  4.50 7.00 7.20 7.50 ;
    END
END OA211X2
MACRO OA211X4
    CLASS CORE ;
    FOREIGN OA211X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  7.10 2.50 7.80 4.20 ;
        RECT  7.50 2.50 7.80 10.55 ;
        RECT  7.25 2.50 7.80 6.30 ;
        RECT  7.50 5.40 7.85 10.55 ;
        RECT  7.15 7.95 7.85 10.55 ;
        RECT  7.50 5.40 8.00 8.45 ;
        RECT  7.15 7.95 8.00 8.45 ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  4.30 5.40 5.35 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 8.05 3.50 11.00 ;
        RECT  4.30 9.55 5.00 11.00 ;
        RECT  0.45 10.70 5.00 11.00 ;
        RECT  5.80 7.95 6.50 11.00 ;
        RECT  8.50 7.95 9.20 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  5.75 2.00 6.45 4.20 ;
        RECT  8.45 2.00 9.15 4.20 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 7.00 1.15 9.55 ;
        RECT  0.55 2.55 1.25 4.00 ;
        RECT  1.90 3.55 2.60 4.25 ;
        RECT  2.10 3.55 2.60 4.95 ;
        RECT  2.10 4.45 3.55 4.95 ;
        RECT  0.55 2.55 3.95 3.05 ;
        RECT  3.05 4.45 3.55 7.50 ;
        RECT  3.25 2.55 3.95 4.00 ;
        RECT  4.30 7.00 5.00 8.55 ;
        RECT  6.35 6.80 7.05 7.50 ;
        RECT  0.45 7.00 7.05 7.50 ;
    END
END OA211X4
MACRO OA21X1
    CLASS CORE ;
    FOREIGN OA21X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.05 1.25 5.05 ;
        RECT  0.75 3.30 1.25 8.80 ;
        RECT  0.75 3.30 1.55 4.05 ;
        RECT  0.75 8.30 2.60 8.80 ;
        RECT  1.90 8.30 2.60 10.00 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.25 8.30 3.95 11.00 ;
        RECT  7.25 8.30 7.95 11.00 ;
        RECT  0.00 11.00 8.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.85 2.00 1.55 2.70 ;
        RECT  5.25 2.00 5.95 3.70 ;
        RECT  0.00 0.00 8.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.95 4.45 2.45 7.80 ;
        RECT  1.95 7.10 2.65 7.80 ;
        RECT  2.55 3.05 3.05 4.95 ;
        RECT  1.95 4.45 3.05 4.95 ;
        RECT  2.55 3.05 3.25 3.75 ;
        RECT  3.90 3.05 4.60 3.75 ;
        RECT  4.10 3.05 4.60 4.65 ;
        RECT  1.95 7.30 5.40 7.80 ;
        RECT  4.90 7.30 5.40 10.00 ;
        RECT  4.90 8.30 5.60 10.00 ;
        RECT  6.60 3.05 7.10 4.65 ;
        RECT  4.10 4.15 7.10 4.65 ;
        RECT  6.60 3.05 7.30 3.75 ;
    END
END OA21X1
MACRO OA21X2
    CLASS CORE ;
    FOREIGN OA21X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.50 3.00 1.00 8.20 ;
        RECT  0.45 3.00 1.15 5.00 ;
        RECT  0.25 4.10 1.15 5.00 ;
        RECT  0.50 7.70 2.75 8.20 ;
        RECT  2.05 7.70 2.75 10.40 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 9.55 1.20 11.00 ;
        RECT  3.40 7.70 4.10 11.00 ;
        RECT  7.25 7.65 7.95 11.00 ;
        RECT  4.90 10.30 7.95 11.00 ;
        RECT  0.00 11.00 8.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 2.70 ;
        RECT  5.90 2.00 6.60 4.00 ;
        RECT  0.00 0.00 8.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.90 6.55 2.60 7.25 ;
        RECT  3.20 3.35 3.70 7.25 ;
        RECT  3.20 3.35 3.90 4.05 ;
        RECT  4.55 3.35 5.25 4.05 ;
        RECT  1.90 6.75 5.40 7.25 ;
        RECT  4.75 3.35 5.25 4.95 ;
        RECT  4.90 6.75 5.40 9.35 ;
        RECT  4.90 7.65 5.60 9.35 ;
        RECT  7.25 3.35 7.75 4.95 ;
        RECT  4.75 4.45 7.75 4.95 ;
        RECT  7.25 3.35 7.95 4.05 ;
    END
END OA21X2
MACRO OA21X4
    CLASS CORE ;
    FOREIGN OA21X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.75 2.55 4.45 ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  2.05 2.75 2.55 7.25 ;
        RECT  2.05 6.75 4.00 7.25 ;
        RECT  3.30 6.75 4.00 10.50 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.55 5.00 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 9.55 1.15 11.00 ;
        RECT  1.95 7.70 2.65 11.00 ;
        RECT  4.65 7.70 5.35 11.00 ;
        RECT  8.65 7.50 9.35 11.00 ;
        RECT  6.15 10.20 9.35 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 4.45 ;
        RECT  3.15 2.00 3.85 4.45 ;
        RECT  5.95 2.00 6.65 3.05 ;
        RECT  8.65 2.00 9.35 3.05 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.00 5.60 3.70 6.30 ;
        RECT  3.00 5.60 5.15 6.10 ;
        RECT  4.65 4.15 5.15 7.25 ;
        RECT  4.65 4.15 5.35 4.85 ;
        RECT  4.65 6.75 6.80 7.25 ;
        RECT  6.00 4.15 6.70 4.85 ;
        RECT  6.30 6.75 6.80 9.20 ;
        RECT  6.30 7.50 7.00 9.20 ;
        RECT  7.30 2.45 7.80 4.65 ;
        RECT  6.00 4.15 7.80 4.65 ;
        RECT  7.30 2.45 8.00 3.15 ;
    END
END OA21X4
MACRO OA221X1
    CLASS CORE ;
    FOREIGN OA221X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.05 3.80 10.40 9.50 ;
        RECT  9.70 7.90 10.40 9.50 ;
        RECT  10.05 3.80 10.55 8.40 ;
        RECT  9.70 7.90 10.55 8.40 ;
        RECT  10.05 3.80 10.95 5.00 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  7.25 6.70 8.15 7.60 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.65 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  0.25 6.70 1.15 7.60 ;
        RECT  4.80 6.75 5.50 7.45 ;
        RECT  0.25 6.95 5.50 7.45 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 9.55 1.20 11.00 ;
        RECT  4.35 8.85 5.05 11.00 ;
        RECT  8.35 8.05 9.05 11.00 ;
        RECT  8.25 10.55 10.75 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.15 2.00 3.85 3.05 ;
        RECT  8.70 2.00 9.40 4.45 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  6.30 8.70 7.40 9.20 ;
        RECT  0.45 2.65 1.15 3.35 ;
        RECT  0.65 2.65 1.15 4.95 ;
        RECT  1.80 2.65 2.50 4.00 ;
        RECT  2.20 7.90 2.70 10.35 ;
        RECT  2.00 8.75 2.70 10.35 ;
        RECT  4.50 2.65 5.20 4.00 ;
        RECT  1.80 3.50 5.20 4.00 ;
        RECT  2.20 7.90 6.80 8.40 ;
        RECT  5.85 2.65 6.35 4.95 ;
        RECT  0.65 4.45 6.35 4.95 ;
        RECT  5.85 2.65 6.55 3.35 ;
        RECT  6.70 5.55 6.80 10.35 ;
        RECT  6.30 5.55 6.80 9.20 ;
        RECT  7.20 2.65 7.90 3.35 ;
        RECT  6.70 8.70 7.40 10.35 ;
        RECT  7.40 2.65 7.90 6.05 ;
        RECT  8.90 5.35 9.60 6.05 ;
        RECT  6.30 5.55 9.60 6.05 ;
    END
END OA221X1
MACRO OA221X2
    CLASS CORE ;
    FOREIGN OA221X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.05 2.80 10.40 10.55 ;
        RECT  9.70 7.15 10.40 10.55 ;
        RECT  10.05 2.80 10.55 7.65 ;
        RECT  9.70 7.15 10.55 7.65 ;
        RECT  10.05 2.80 10.75 5.00 ;
        RECT  10.05 3.80 10.95 5.00 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  7.25 6.70 8.15 7.60 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.65 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  0.25 6.70 1.15 7.60 ;
        RECT  4.80 6.75 5.50 7.45 ;
        RECT  0.25 6.95 5.50 7.45 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 9.55 1.20 11.00 ;
        RECT  4.35 8.85 5.05 11.00 ;
        RECT  8.35 8.05 9.05 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.15 2.00 3.85 3.05 ;
        RECT  8.70 2.00 9.40 4.45 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  6.30 8.70 7.40 9.20 ;
        RECT  0.45 2.65 1.15 3.35 ;
        RECT  0.65 2.65 1.15 4.95 ;
        RECT  1.80 2.65 2.50 4.00 ;
        RECT  2.20 7.90 2.70 10.35 ;
        RECT  2.00 8.75 2.70 10.35 ;
        RECT  4.50 2.65 5.20 4.00 ;
        RECT  1.80 3.50 5.20 4.00 ;
        RECT  2.20 7.90 6.80 8.40 ;
        RECT  5.85 2.65 6.35 4.95 ;
        RECT  0.65 4.45 6.35 4.95 ;
        RECT  5.85 2.65 6.55 3.35 ;
        RECT  6.70 5.55 6.80 10.35 ;
        RECT  6.30 5.55 6.80 9.20 ;
        RECT  7.20 2.65 7.90 3.35 ;
        RECT  6.70 8.70 7.40 10.35 ;
        RECT  7.40 2.65 7.90 6.05 ;
        RECT  8.90 5.35 9.60 6.05 ;
        RECT  6.30 5.55 9.60 6.05 ;
    END
END OA221X2
MACRO OA221X4
    CLASS CORE ;
    FOREIGN OA221X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.05 2.80 10.55 10.55 ;
        RECT  9.95 7.15 10.65 10.55 ;
        RECT  10.05 2.80 10.75 5.00 ;
        RECT  10.05 4.10 10.95 5.00 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  7.25 6.70 8.15 7.60 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.65 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        RECT  0.65 5.40 1.15 7.25 ;
        RECT  0.65 6.75 5.75 7.25 ;
        RECT  5.05 6.75 5.75 7.45 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.55 9.55 1.25 11.00 ;
        RECT  4.60 8.85 5.30 11.00 ;
        RECT  8.60 7.20 9.30 11.00 ;
        RECT  11.30 7.20 12.00 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.15 2.00 3.85 3.05 ;
        RECT  8.70 2.00 9.40 4.45 ;
        RECT  11.40 2.00 12.10 4.45 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 2.65 1.15 3.35 ;
        RECT  0.65 2.65 1.15 4.95 ;
        RECT  1.80 2.65 2.50 4.00 ;
        RECT  2.45 7.90 2.95 10.35 ;
        RECT  2.25 8.75 2.95 10.35 ;
        RECT  4.50 2.65 5.20 4.00 ;
        RECT  1.80 3.50 5.20 4.00 ;
        RECT  2.45 7.90 6.80 8.40 ;
        RECT  5.85 2.65 6.35 4.95 ;
        RECT  0.65 4.45 6.35 4.95 ;
        RECT  5.85 2.65 6.55 3.35 ;
        RECT  6.30 5.55 6.80 9.20 ;
        RECT  6.30 8.70 7.65 9.20 ;
        RECT  7.20 2.65 7.90 3.35 ;
        RECT  6.95 8.70 7.65 10.35 ;
        RECT  7.40 2.65 7.90 6.05 ;
        RECT  8.90 5.35 9.60 6.05 ;
        RECT  6.30 5.55 9.60 6.05 ;
    END
END OA221X4
MACRO OA222X1
    CLASS CORE ;
    FOREIGN OA222X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.40 8.85 11.15 10.45 ;
        RECT  11.45 3.75 12.00 9.35 ;
        RECT  10.40 8.85 12.00 9.35 ;
        RECT  11.45 3.75 12.15 6.30 ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  8.65 6.70 9.55 7.60 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  7.25 6.70 8.15 7.60 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        RECT  0.65 5.40 1.15 7.25 ;
        RECT  0.65 6.75 5.50 7.25 ;
        RECT  4.80 6.75 5.50 7.45 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 9.60 1.15 11.00 ;
        RECT  4.35 8.85 5.05 11.00 ;
        RECT  9.05 8.75 9.75 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.15 2.00 3.85 3.05 ;
        RECT  10.10 2.00 10.80 4.45 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  6.30 8.75 7.40 9.25 ;
        RECT  0.45 2.65 1.15 3.35 ;
        RECT  0.65 2.65 1.15 4.95 ;
        RECT  1.80 2.65 2.50 4.00 ;
        RECT  2.20 7.90 2.70 10.35 ;
        RECT  2.00 8.75 2.70 10.35 ;
        RECT  4.50 2.65 5.20 4.00 ;
        RECT  1.80 3.50 5.20 4.00 ;
        RECT  2.20 7.90 6.80 8.40 ;
        RECT  5.85 2.45 6.35 4.95 ;
        RECT  0.65 4.45 6.35 4.95 ;
        RECT  5.85 2.45 6.55 3.65 ;
        RECT  6.70 5.55 6.80 10.35 ;
        RECT  6.30 5.55 6.80 9.25 ;
        RECT  6.70 8.75 7.40 10.35 ;
        RECT  7.20 3.40 7.70 6.05 ;
        RECT  7.20 3.40 7.90 4.10 ;
        RECT  5.85 2.45 9.25 2.95 ;
        RECT  8.55 2.45 9.25 3.65 ;
        RECT  9.95 5.35 10.65 6.05 ;
        RECT  6.30 5.55 10.65 6.05 ;
    END
END OA222X1
MACRO OA222X2
    CLASS CORE ;
    FOREIGN OA222X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.55 7.85 11.30 10.55 ;
        RECT  11.45 2.75 12.00 8.35 ;
        RECT  10.55 7.85 12.00 8.35 ;
        RECT  11.45 2.75 12.15 6.30 ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  8.65 6.70 9.55 7.60 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  7.25 6.70 8.15 7.60 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        RECT  0.65 5.40 1.15 7.25 ;
        RECT  0.65 6.75 5.50 7.25 ;
        RECT  4.80 6.75 5.50 7.45 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 9.60 1.15 11.00 ;
        RECT  4.35 8.85 5.05 11.00 ;
        RECT  9.20 8.05 9.90 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.15 2.00 3.85 3.05 ;
        RECT  10.10 2.00 10.80 4.45 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  6.30 8.75 7.40 9.25 ;
        RECT  0.45 2.65 1.15 3.35 ;
        RECT  0.65 2.65 1.15 4.95 ;
        RECT  1.80 2.65 2.50 4.00 ;
        RECT  2.20 7.90 2.70 10.35 ;
        RECT  2.00 8.75 2.70 10.35 ;
        RECT  4.50 2.65 5.20 4.00 ;
        RECT  1.80 3.50 5.20 4.00 ;
        RECT  2.20 7.90 6.80 8.40 ;
        RECT  5.85 2.45 6.35 4.95 ;
        RECT  0.65 4.45 6.35 4.95 ;
        RECT  5.85 2.45 6.55 3.65 ;
        RECT  6.70 5.55 6.80 10.35 ;
        RECT  6.30 5.55 6.80 9.25 ;
        RECT  6.70 8.75 7.40 10.35 ;
        RECT  7.20 3.40 7.70 6.05 ;
        RECT  7.20 3.40 7.90 4.10 ;
        RECT  5.85 2.45 9.25 2.95 ;
        RECT  8.55 2.45 9.25 3.65 ;
        RECT  10.10 5.35 10.80 6.05 ;
        RECT  6.30 5.55 10.80 6.05 ;
    END
END OA222X2
MACRO OA222X4
    CLASS CORE ;
    FOREIGN OA222X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.75 6.50 11.25 10.55 ;
        RECT  10.55 7.85 11.25 10.55 ;
        RECT  11.45 2.75 12.00 7.00 ;
        RECT  10.75 6.50 12.00 7.00 ;
        RECT  11.45 2.75 12.15 6.30 ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  8.65 6.70 9.55 7.60 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  7.25 6.70 8.15 7.60 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        RECT  0.65 5.40 1.15 7.25 ;
        RECT  0.65 6.75 5.50 7.25 ;
        RECT  4.80 6.75 5.50 7.45 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 9.55 1.15 11.00 ;
        RECT  4.35 8.85 5.05 11.00 ;
        RECT  9.20 8.05 9.90 11.00 ;
        RECT  11.90 8.05 12.60 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.15 2.00 3.85 3.05 ;
        RECT  10.10 2.00 10.80 4.45 ;
        RECT  12.80 2.00 13.50 4.45 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  6.30 8.75 7.40 9.25 ;
        RECT  0.45 2.65 1.15 3.35 ;
        RECT  0.65 2.65 1.15 4.95 ;
        RECT  1.80 2.65 2.50 4.00 ;
        RECT  2.20 7.90 2.70 10.35 ;
        RECT  2.00 8.75 2.70 10.35 ;
        RECT  4.50 2.65 5.20 4.00 ;
        RECT  1.80 3.50 5.20 4.00 ;
        RECT  2.20 7.90 6.80 8.40 ;
        RECT  5.85 2.45 6.35 4.95 ;
        RECT  0.65 4.45 6.35 4.95 ;
        RECT  5.85 2.45 6.55 3.65 ;
        RECT  6.70 5.55 6.80 10.35 ;
        RECT  6.30 5.55 6.80 9.25 ;
        RECT  6.70 8.75 7.40 10.35 ;
        RECT  7.20 3.40 7.70 6.05 ;
        RECT  7.20 3.40 7.90 4.10 ;
        RECT  5.85 2.45 9.25 2.95 ;
        RECT  8.55 2.45 9.25 3.65 ;
        RECT  10.30 5.35 11.00 6.05 ;
        RECT  6.30 5.55 11.00 6.05 ;
    END
END OA222X4
MACRO OA22X1
    CLASS CORE ;
    FOREIGN OA22X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.25 3.60 0.75 10.25 ;
        RECT  0.25 9.75 1.70 10.25 ;
        RECT  0.25 3.60 1.25 5.00 ;
        RECT  0.25 3.60 1.65 4.30 ;
        RECT  1.00 9.75 1.70 10.45 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 6.70 8.15 7.60 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.75 5.35 6.75 6.35 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.60 6.70 2.55 7.60 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 8.00 5.35 8.90 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.35 9.35 3.05 11.00 ;
        RECT  7.25 9.30 7.95 11.00 ;
        RECT  0.00 11.00 8.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 2.00 1.65 2.80 ;
        RECT  3.25 2.00 3.95 2.50 ;
        RECT  6.65 2.00 7.35 2.80 ;
        RECT  0.00 0.00 8.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.45 8.05 2.15 8.75 ;
        RECT  2.25 3.35 2.75 6.25 ;
        RECT  2.25 5.75 3.95 6.25 ;
        RECT  1.45 8.05 4.00 8.55 ;
        RECT  3.25 3.15 3.95 3.85 ;
        RECT  3.25 4.55 3.95 5.25 ;
        RECT  3.25 5.75 3.95 6.60 ;
        RECT  3.50 7.05 4.00 10.25 ;
        RECT  3.25 4.75 4.95 5.25 ;
        RECT  3.50 9.75 5.60 10.25 ;
        RECT  4.45 4.75 4.95 7.55 ;
        RECT  3.50 7.05 4.95 7.55 ;
        RECT  4.90 9.75 5.60 10.45 ;
        RECT  2.25 3.35 7.35 3.85 ;
        RECT  6.65 3.35 7.35 4.15 ;
    END
END OA22X1
MACRO OA22X2
    CLASS CORE ;
    FOREIGN OA22X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.45 1.15 4.05 ;
        RECT  0.25 5.40 1.15 6.30 ;
        RECT  0.65 2.45 1.15 10.55 ;
        RECT  0.50 9.85 2.10 10.55 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 4.10 8.15 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 6.70 6.75 7.60 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.55 7.60 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 8.00 5.35 8.90 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  7.25 9.30 7.95 11.00 ;
        RECT  0.00 11.00 8.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 3.85 ;
        RECT  3.90 2.00 4.60 2.25 ;
        RECT  0.00 0.00 8.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.85 8.05 3.50 8.75 ;
        RECT  3.00 4.50 3.50 9.85 ;
        RECT  3.85 4.30 4.55 5.00 ;
        RECT  3.00 4.50 4.55 5.00 ;
        RECT  3.95 5.65 4.65 6.35 ;
        RECT  3.00 9.35 5.60 9.85 ;
        RECT  3.90 2.90 5.50 3.60 ;
        RECT  5.00 2.90 5.50 6.15 ;
        RECT  3.95 5.65 5.50 6.15 ;
        RECT  4.90 9.35 5.60 10.45 ;
        RECT  6.70 2.65 7.40 3.40 ;
        RECT  3.90 2.90 7.40 3.40 ;
    END
END OA22X2
MACRO OA22X4
    CLASS CORE ;
    FOREIGN OA22X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  2.20 8.05 3.05 8.55 ;
        RECT  1.90 2.45 2.70 4.50 ;
        RECT  1.65 5.40 2.70 6.30 ;
        RECT  2.35 2.45 2.70 10.55 ;
        RECT  2.20 2.45 2.70 8.55 ;
        RECT  2.35 8.05 3.05 10.55 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.55 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.35 7.60 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.80 6.70 6.75 7.60 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.00 8.10 1.70 11.00 ;
        RECT  3.70 9.00 4.40 11.00 ;
        RECT  8.55 7.90 9.25 11.00 ;
        RECT  5.20 10.55 9.35 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.55 2.00 1.25 4.50 ;
        RECT  3.55 2.00 5.15 3.05 ;
        RECT  5.95 2.00 6.65 3.05 ;
        RECT  8.65 2.00 9.35 3.05 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.15 5.65 4.00 6.35 ;
        RECT  3.50 5.65 4.00 8.55 ;
        RECT  3.50 3.50 4.20 5.05 ;
        RECT  4.85 4.45 5.35 6.15 ;
        RECT  3.15 5.65 5.35 6.15 ;
        RECT  4.85 4.45 5.55 5.15 ;
        RECT  3.50 8.05 6.90 8.55 ;
        RECT  6.20 3.50 6.90 5.05 ;
        RECT  6.20 8.05 6.90 9.65 ;
        RECT  7.30 2.45 7.80 4.00 ;
        RECT  3.50 3.50 7.80 4.00 ;
        RECT  7.30 2.45 8.00 3.15 ;
    END
END OA22X4
MACRO OA311X1
    CLASS CORE ;
    FOREIGN OA311X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.35 6.40 8.85 9.30 ;
        RECT  8.15 7.70 8.85 9.30 ;
        RECT  9.70 3.75 10.45 4.45 ;
        RECT  9.95 3.75 10.45 6.90 ;
        RECT  8.35 6.40 10.45 6.90 ;
        RECT  9.95 5.40 10.95 6.30 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.80 7.70 4.50 11.00 ;
        RECT  5.30 10.10 6.00 11.00 ;
        RECT  6.80 7.70 7.50 11.00 ;
        RECT  10.05 9.55 10.75 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.75 ;
        RECT  3.15 2.00 3.85 3.75 ;
        RECT  8.35 2.00 9.05 4.45 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 6.75 1.15 10.05 ;
        RECT  1.75 3.30 2.50 4.75 ;
        RECT  4.50 3.30 5.20 4.75 ;
        RECT  1.75 4.25 5.20 4.75 ;
        RECT  5.30 6.75 6.00 8.40 ;
        RECT  6.85 3.30 7.70 4.00 ;
        RECT  7.20 3.30 7.70 7.25 ;
        RECT  0.45 6.75 7.70 7.25 ;
        RECT  7.20 5.25 9.50 5.75 ;
        RECT  8.80 5.25 9.50 5.95 ;
    END
END OA311X1
MACRO OA311X2
    CLASS CORE ;
    FOREIGN OA311X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.35 6.40 8.85 10.50 ;
        RECT  8.15 7.70 8.85 10.50 ;
        RECT  9.70 2.75 10.45 4.45 ;
        RECT  9.95 2.75 10.45 6.90 ;
        RECT  8.35 6.40 10.45 6.90 ;
        RECT  9.95 5.40 10.95 6.30 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.80 7.70 4.50 11.00 ;
        RECT  5.30 10.10 6.00 11.00 ;
        RECT  6.80 7.70 7.50 11.00 ;
        RECT  9.85 9.55 10.55 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.75 ;
        RECT  3.15 2.00 3.85 3.75 ;
        RECT  8.35 2.00 9.05 4.45 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 6.75 1.15 10.05 ;
        RECT  1.75 3.30 2.50 4.75 ;
        RECT  4.50 3.30 5.20 4.75 ;
        RECT  1.75 4.25 5.20 4.75 ;
        RECT  5.30 6.75 6.00 8.40 ;
        RECT  6.85 3.30 7.70 4.00 ;
        RECT  7.20 3.30 7.70 7.25 ;
        RECT  0.45 6.75 7.70 7.25 ;
        RECT  7.20 5.25 9.50 5.75 ;
        RECT  8.80 5.25 9.50 5.95 ;
    END
END OA311X2
MACRO OA311X4
    CLASS CORE ;
    FOREIGN OA311X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.35 6.00 8.85 10.50 ;
        RECT  8.15 7.70 8.85 10.50 ;
        RECT  9.70 2.45 10.45 4.35 ;
        RECT  9.95 2.45 10.45 6.50 ;
        RECT  9.95 5.40 10.95 6.50 ;
        RECT  8.35 6.00 10.95 6.50 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.80 7.70 4.50 11.00 ;
        RECT  5.30 10.10 6.00 11.00 ;
        RECT  6.80 7.70 7.50 11.00 ;
        RECT  9.50 7.70 10.20 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.75 ;
        RECT  3.15 2.00 3.85 3.75 ;
        RECT  8.35 2.00 9.05 4.35 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 6.75 1.15 10.05 ;
        RECT  1.75 3.30 2.50 4.75 ;
        RECT  4.50 3.30 5.20 4.75 ;
        RECT  1.75 4.25 5.20 4.75 ;
        RECT  5.30 6.75 6.00 8.40 ;
        RECT  6.85 3.30 7.70 4.00 ;
        RECT  7.20 3.30 7.70 7.25 ;
        RECT  0.45 6.75 7.70 7.25 ;
        RECT  7.20 4.85 9.50 5.35 ;
        RECT  8.80 4.85 9.50 5.55 ;
    END
END OA311X4
MACRO OA31X1
    CLASS CORE ;
    FOREIGN OA31X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.75 3.35 0.90 9.40 ;
        RECT  0.40 8.90 1.60 9.40 ;
        RECT  0.40 4.05 0.90 9.40 ;
        RECT  0.75 3.35 1.25 5.05 ;
        RECT  0.25 4.05 1.25 5.05 ;
        RECT  0.90 8.90 1.60 10.50 ;
        RECT  0.75 3.35 1.75 4.05 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.35 7.60 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  5.85 6.70 6.75 7.60 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.25 9.00 2.95 11.00 ;
        RECT  7.25 8.85 7.95 11.00 ;
        RECT  0.00 11.00 8.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.05 2.00 1.75 2.60 ;
        RECT  3.00 2.00 3.70 3.45 ;
        RECT  4.55 2.00 5.25 3.20 ;
        RECT  7.25 2.00 7.95 3.25 ;
        RECT  0.00 0.00 8.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.35 8.05 4.60 8.25 ;
        RECT  1.35 7.75 2.05 8.45 ;
        RECT  3.00 5.45 3.70 6.15 ;
        RECT  3.00 4.10 3.70 4.80 ;
        RECT  3.20 5.45 3.70 8.55 ;
        RECT  1.35 7.75 3.70 8.25 ;
        RECT  3.20 8.05 4.60 8.55 ;
        RECT  3.90 8.05 4.60 10.45 ;
        RECT  5.90 2.55 6.40 4.60 ;
        RECT  3.00 4.10 6.40 4.60 ;
        RECT  5.90 2.55 6.60 3.25 ;
    END
END OA31X1
#MACRO OA31X2
#    CLASS CORE ;
#    FOREIGN OA31X2 0.00 0.00  ;
#    ORIGIN 0.00 0.00 ;
#    SIZE 9.80 BY 13.00 ;
#    SYMMETRY x y r90 ;
#    SITE core ;
#    PIN Q
#        DIRECTION OUTPUT ;
#        ANTENNADIFFAREA 1.0 ;
#        PORT
#        LAYER M1M ;
#        RECT  1.65 4.10 2.80 5.00 ;
#        RECT  2.30 2.80 2.50 10.55 ;
#        RECT  1.80 2.80 2.50 5.00 ;
#        RECT  2.30 4.10 2.80 10.55 ;
#        RECT  2.30 8.95 3.00 10.55 ;
#        END
#    END Q
#    PIN D
#        DIRECTION INPUT ;
#        ANTENNAGATEAREA 0.70 ;
#        PORT
#        LAYER M1M ;
#        RECT  4.45 6.70 5.35 7.60 ;
#        END
#    END D
#    PIN C
#        DIRECTION INPUT ;
#        ANTENNAGATEAREA 1.40 ;
#        PORT
#        LAYER M1M ;
#        RECT  5.85 5.40 6.75 6.30 ;
#        END
#    END C
#    PIN B
#        DIRECTION INPUT ;
#        ANTENNAGATEAREA 1.40 ;
#        PORT
#        LAYER M1M ;
#        RECT  7.25 6.70 8.15 7.60 ;
#        END
#    END B
#    PIN A
#        DIRECTION INPUT ;
#        ANTENNAGATEAREA 1.40 ;
#        PORT
#        LAYER M1M ;
#        RECT  8.65 5.40 9.55 6.30 ;
#        END
#    END A
#    PIN vdd!
#        DIRECTION INOUT ;
#        USE power ;
#        SHAPE ABUTMENT ;
#        PORT
#        LAYER M1M ;
#        RECT  0.95 9.00 1.65 11.00 ;
#        RECT  3.65 9.00 4.35 11.00 ;
#        RECT  8.65 8.85 9.35 11.00 ;
#        RECT  0.00 11.00 9.80 13.00 ;
#        END
#    END vdd!
#    PIN gnd!
#        DIRECTION INOUT ;
#        USE ground ;
#        SHAPE ABUTMENT ;
#        PORT
#        LAYER M1M ;
#        RECT  0.45 2.00 1.15 4.40 ;
#        RECT  5.95 2.00 6.65 3.20 ;
#        RECT  8.65 2.00 9.35 3.25 ;
#        RECT  0.00 0.00 9.80 2.00 ;
#        END
#    END gnd!
#    OBS
#        LAYER M1M ;
#        RECT  3.45 4.35 3.95 8.55 ;
#        RECT  3.25 7.75 3.95 8.55 ;
#        RECT  3.45 4.35 4.15 5.05 ;
#        RECT  4.60 2.55 5.30 3.25 ;
#        RECT  3.25 8.05 6.00 8.55 ;
#        RECT  4.80 2.55 5.30 5.05 ;
#        RECT  4.80 4.35 5.50 5.05 ;
#        RECT  5.30 8.05 6.00 10.45 ;
#        RECT  7.30 2.55 7.80 4.85 ;
#        RECT  4.80 4.35 7.80 4.85 ;
#        RECT  7.30 2.55 8.00 3.25 ;
#    END
#END OA31X2
MACRO OA31X4
    CLASS CORE ;
    FOREIGN OA31X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.65 4.10 2.80 5.00 ;
        RECT  2.30 2.55 2.50 10.55 ;
        RECT  1.80 2.55 2.50 5.00 ;
        RECT  2.30 4.10 2.80 10.55 ;
        RECT  2.30 7.75 3.00 10.55 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.70 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.55 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.95 7.75 1.65 11.00 ;
        RECT  3.65 7.75 4.35 11.00 ;
        RECT  8.65 7.70 9.35 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 4.40 ;
        RECT  5.95 2.00 6.65 3.20 ;
        RECT  8.65 2.00 9.35 3.25 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.45 4.30 3.95 7.30 ;
        RECT  3.25 6.60 3.95 7.30 ;
        RECT  3.45 4.30 4.15 5.00 ;
        RECT  4.60 2.55 5.30 3.25 ;
        RECT  3.25 6.80 6.00 7.30 ;
        RECT  4.80 2.55 5.30 4.95 ;
        RECT  4.80 4.25 5.50 4.95 ;
        RECT  5.30 6.80 6.00 10.40 ;
        RECT  7.30 2.55 7.80 4.75 ;
        RECT  4.80 4.25 7.80 4.75 ;
        RECT  7.30 2.55 8.00 3.25 ;
    END
END OA31X4
MACRO OA321X1
    CLASS CORE ;
    FOREIGN OA321X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  9.75 2.45 10.45 3.15 ;
        RECT  9.35 8.85 10.05 10.45 ;
        RECT  10.05 2.45 10.45 9.35 ;
        RECT  9.95 2.45 10.45 5.00 ;
        RECT  10.05 4.10 10.55 9.35 ;
        RECT  9.35 8.85 10.55 9.35 ;
        RECT  9.95 4.10 10.95 5.00 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  8.65 6.70 9.55 7.60 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  5.85 6.70 6.75 7.60 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.35 7.60 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.65 2.85 7.60 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 4.05 5.05 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.80 8.50 4.50 11.00 ;
        RECT  8.00 9.00 8.70 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 2.75 ;
        RECT  3.15 2.00 3.85 2.70 ;
        RECT  8.30 2.00 9.00 3.00 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.65 5.65 1.15 10.45 ;
        RECT  0.45 8.65 1.15 10.45 ;
        RECT  1.80 2.55 2.50 3.65 ;
        RECT  4.50 2.55 5.20 3.65 ;
        RECT  1.80 3.15 5.20 3.65 ;
        RECT  4.70 2.55 5.20 5.15 ;
        RECT  4.70 4.45 6.15 5.15 ;
        RECT  5.85 2.45 7.30 3.15 ;
        RECT  6.30 8.05 7.00 10.45 ;
        RECT  6.80 2.45 7.30 5.15 ;
        RECT  6.80 4.45 7.50 5.15 ;
        RECT  7.20 5.65 7.70 8.55 ;
        RECT  6.30 8.05 7.70 8.55 ;
        RECT  8.15 3.85 8.85 4.55 ;
        RECT  8.35 3.85 8.85 6.15 ;
        RECT  8.35 5.45 9.55 6.15 ;
        RECT  0.65 5.65 9.55 6.15 ;
    END
END OA321X1
MACRO OA321X2
    CLASS CORE ;
    FOREIGN OA321X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  9.75 2.45 10.45 3.15 ;
        RECT  9.35 8.80 10.05 10.45 ;
        RECT  10.05 2.45 10.45 9.35 ;
        RECT  9.95 2.45 10.45 5.00 ;
        RECT  10.05 4.10 10.55 9.35 ;
        RECT  9.35 8.80 10.55 9.35 ;
        RECT  9.95 4.10 10.95 5.00 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  8.65 6.70 9.55 7.60 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  5.85 6.70 6.75 7.60 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.35 7.60 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.55 2.80 7.60 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 4.05 5.05 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.80 8.50 4.50 11.00 ;
        RECT  8.00 9.00 8.70 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 2.75 ;
        RECT  3.15 2.00 3.85 2.70 ;
        RECT  8.30 2.00 9.00 3.00 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.65 5.60 1.15 10.45 ;
        RECT  0.45 8.65 1.15 10.45 ;
        RECT  1.80 2.55 2.50 3.65 ;
        RECT  4.50 2.55 5.20 3.65 ;
        RECT  1.80 3.15 5.20 3.65 ;
        RECT  4.70 2.55 5.20 5.15 ;
        RECT  4.70 4.45 6.15 5.15 ;
        RECT  5.85 2.45 7.30 3.15 ;
        RECT  6.30 8.05 7.00 10.45 ;
        RECT  6.80 2.45 7.30 5.15 ;
        RECT  6.80 4.45 7.50 5.15 ;
        RECT  7.20 5.60 7.70 8.55 ;
        RECT  6.30 8.05 7.70 8.55 ;
        RECT  8.15 3.85 8.85 4.55 ;
        RECT  8.35 3.85 8.85 6.10 ;
        RECT  8.35 5.40 9.55 6.10 ;
        RECT  0.65 5.60 9.55 6.10 ;
    END
END OA321X2
MACRO OA321X4
    CLASS CORE ;
    FOREIGN OA321X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.00 7.10 10.30 10.55 ;
        RECT  9.60 8.80 10.30 10.55 ;
        RECT  10.00 7.10 10.50 9.35 ;
        RECT  9.60 8.80 10.50 9.35 ;
        RECT  11.30 2.45 12.00 4.35 ;
        RECT  11.45 2.45 12.00 7.60 ;
        RECT  11.45 6.70 12.35 7.60 ;
        RECT  10.00 7.10 12.35 7.60 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  8.65 6.50 9.55 7.60 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  5.85 6.70 6.75 7.60 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.35 7.60 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 4.30 5.05 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  4.10 8.35 4.80 11.00 ;
        RECT  8.25 8.40 8.95 11.00 ;
        RECT  10.95 8.40 11.65 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 2.75 ;
        RECT  3.15 2.00 3.85 2.70 ;
        RECT  7.40 2.00 9.15 2.90 ;
        RECT  9.95 2.00 10.65 4.50 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.95 6.90 1.45 10.45 ;
        RECT  0.75 8.65 1.45 10.45 ;
        RECT  1.80 2.55 2.50 3.65 ;
        RECT  3.10 5.50 3.60 7.40 ;
        RECT  0.95 6.90 3.60 7.40 ;
        RECT  4.50 2.55 5.25 3.65 ;
        RECT  1.80 3.15 5.25 3.65 ;
        RECT  4.75 2.55 5.25 5.05 ;
        RECT  4.75 4.35 6.45 5.05 ;
        RECT  5.85 2.45 6.55 3.85 ;
        RECT  5.85 3.35 7.80 3.85 ;
        RECT  7.20 5.50 7.30 10.00 ;
        RECT  6.60 8.20 7.30 10.00 ;
        RECT  7.20 5.50 7.70 8.70 ;
        RECT  6.60 8.20 7.70 8.70 ;
        RECT  7.10 3.35 7.80 5.05 ;
        RECT  8.45 4.35 9.15 6.00 ;
        RECT  10.30 5.30 11.00 6.00 ;
        RECT  3.10 5.50 11.00 6.00 ;
    END
END OA321X4
MACRO OA322X1
    CLASS CORE ;
    FOREIGN OA322X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.20 8.95 10.90 10.55 ;
        RECT  11.45 3.70 11.95 9.50 ;
        RECT  10.20 8.95 11.95 9.50 ;
        RECT  11.45 3.70 12.15 4.40 ;
        RECT  11.45 6.70 12.35 7.60 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  8.15 6.30 9.55 7.00 ;
        RECT  8.65 6.30 9.55 7.60 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  10.05 6.65 10.95 7.60 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  5.85 6.70 6.75 7.60 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.35 7.60 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.60 2.85 7.60 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 4.10 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.80 8.25 4.50 11.00 ;
        RECT  8.70 8.20 9.55 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 2.75 ;
        RECT  3.15 2.00 3.85 2.70 ;
        RECT  10.10 2.00 10.80 4.40 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.65 5.65 1.15 10.45 ;
        RECT  0.45 8.65 1.15 10.45 ;
        RECT  1.80 2.55 2.50 3.65 ;
        RECT  4.50 2.55 5.20 3.65 ;
        RECT  1.80 3.15 5.20 3.65 ;
        RECT  4.70 2.55 5.20 5.00 ;
        RECT  4.70 4.50 6.15 5.00 ;
        RECT  5.45 4.50 6.15 5.20 ;
        RECT  5.85 2.55 7.15 3.25 ;
        RECT  6.35 8.30 7.05 9.90 ;
        RECT  6.65 2.55 7.15 4.90 ;
        RECT  0.65 5.65 7.70 6.15 ;
        RECT  6.65 4.20 7.65 4.90 ;
        RECT  7.20 5.35 7.70 8.80 ;
        RECT  6.35 8.30 7.70 8.80 ;
        RECT  7.60 2.55 8.65 3.25 ;
        RECT  7.20 5.35 8.65 5.85 ;
        RECT  8.15 2.55 8.65 5.85 ;
        RECT  0.65 5.65 8.65 5.85 ;
        RECT  8.15 4.80 9.10 5.55 ;
        RECT  8.15 5.05 11.00 5.55 ;
        RECT  10.30 4.85 11.00 5.55 ;
        RECT  7.20 5.35 11.00 5.55 ;
    END
END OA322X1
MACRO OA322X2
    CLASS CORE ;
    FOREIGN OA322X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.45 2.70 11.95 10.55 ;
        RECT  10.20 8.95 11.95 10.55 ;
        RECT  11.45 2.70 12.15 4.40 ;
        RECT  11.45 6.70 12.35 7.60 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  8.15 6.30 9.55 7.00 ;
        RECT  8.65 6.30 9.55 7.60 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  10.05 6.65 10.95 7.60 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  5.85 6.70 6.75 7.60 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.35 7.60 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.60 2.85 7.60 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 4.10 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.80 8.25 4.50 11.00 ;
        RECT  8.70 8.20 9.55 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 2.75 ;
        RECT  3.15 2.00 3.85 2.70 ;
        RECT  10.10 2.00 10.80 4.40 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.65 5.65 1.15 10.45 ;
        RECT  0.45 8.65 1.15 10.45 ;
        RECT  1.80 2.55 2.50 3.65 ;
        RECT  4.55 2.55 5.25 3.65 ;
        RECT  1.80 3.15 5.25 3.65 ;
        RECT  4.75 2.55 5.25 5.00 ;
        RECT  4.75 4.50 6.15 5.00 ;
        RECT  5.45 4.50 6.15 5.20 ;
        RECT  5.95 2.55 7.15 3.25 ;
        RECT  6.35 8.30 7.05 9.90 ;
        RECT  6.65 2.55 7.15 4.90 ;
        RECT  0.65 5.65 7.70 6.15 ;
        RECT  6.65 4.20 7.65 4.90 ;
        RECT  7.20 5.35 7.70 8.80 ;
        RECT  6.35 8.30 7.70 8.80 ;
        RECT  7.60 2.55 8.65 3.25 ;
        RECT  7.20 5.35 8.65 5.85 ;
        RECT  8.15 2.55 8.65 5.85 ;
        RECT  0.65 5.65 8.65 5.85 ;
        RECT  8.15 4.85 9.10 5.55 ;
        RECT  8.15 5.05 11.00 5.55 ;
        RECT  10.30 4.85 11.00 5.55 ;
        RECT  7.20 5.35 11.00 5.55 ;
    END
END OA322X2
MACRO OA322X4
    CLASS CORE ;
    FOREIGN OA322X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.45 2.70 12.15 4.40 ;
        RECT  11.65 2.70 12.15 10.55 ;
        RECT  11.45 8.95 12.15 10.55 ;
        RECT  11.45 6.70 12.35 7.60 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.60 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  9.75 5.35 10.95 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.60 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.40 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  1.65 5.55 2.90 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 3.95 5.00 ;
        RECT  3.05 4.10 4.30 4.85 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  4.35 8.30 5.05 11.00 ;
        RECT  9.20 8.30 10.80 11.00 ;
        RECT  12.80 8.30 13.50 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 2.75 ;
        RECT  3.15 2.00 3.85 2.70 ;
        RECT  10.10 2.00 10.80 4.40 ;
        RECT  12.80 2.00 13.50 4.40 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  8.40 4.25 9.10 4.95 ;
        RECT  1.00 7.35 1.70 10.20 ;
        RECT  1.80 2.55 2.50 3.65 ;
        RECT  4.50 2.55 5.25 3.65 ;
        RECT  1.80 3.15 5.25 3.65 ;
        RECT  4.75 2.55 5.25 4.95 ;
        RECT  4.75 4.25 6.15 4.95 ;
        RECT  5.95 2.55 7.15 3.25 ;
        RECT  6.65 2.55 7.15 4.95 ;
        RECT  6.85 7.35 7.55 9.90 ;
        RECT  6.65 4.25 7.65 4.95 ;
        RECT  7.60 2.55 8.90 3.25 ;
        RECT  8.60 2.55 8.90 7.85 ;
        RECT  8.40 2.55 8.90 4.95 ;
        RECT  8.60 4.25 9.10 7.85 ;
        RECT  10.30 7.15 11.00 7.85 ;
        RECT  1.00 7.35 11.00 7.85 ;
    END
END OA322X4
MACRO OA32X1
    CLASS CORE ;
    FOREIGN OA32X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.15 3.75 9.55 4.45 ;
        RECT  8.65 3.75 9.15 10.45 ;
        RECT  7.65 9.75 9.15 10.45 ;
        RECT  8.65 3.75 9.55 5.00 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.35 7.60 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 6.70 8.15 7.60 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 8.30 1.15 11.00 ;
        RECT  6.30 9.30 7.00 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.10 ;
        RECT  3.15 2.00 3.85 3.10 ;
        RECT  8.15 2.00 8.85 2.95 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 2.45 2.55 3.15 ;
        RECT  2.05 2.45 2.55 4.25 ;
        RECT  3.80 8.15 4.50 10.45 ;
        RECT  4.50 2.45 4.70 5.60 ;
        RECT  4.00 3.75 4.70 5.60 ;
        RECT  4.50 2.45 5.00 4.25 ;
        RECT  2.05 3.75 5.00 4.25 ;
        RECT  4.50 2.45 5.20 3.15 ;
        RECT  5.35 4.85 6.30 5.55 ;
        RECT  5.80 2.45 6.30 8.65 ;
        RECT  5.80 2.45 6.55 3.15 ;
        RECT  3.80 8.15 7.95 8.65 ;
        RECT  7.25 8.15 7.95 8.85 ;
        RECT  7.45 5.45 8.15 6.15 ;
        RECT  5.80 5.65 8.15 6.15 ;
    END
END OA32X1
MACRO OA32X2
    CLASS CORE ;
    FOREIGN OA32X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.15 6.70 8.65 10.55 ;
        RECT  7.95 8.95 8.65 10.55 ;
        RECT  8.80 2.75 9.55 4.35 ;
        RECT  9.05 2.75 9.55 7.60 ;
        RECT  8.15 6.70 9.55 7.60 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.35 7.60 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 6.70 6.75 7.60 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.55 8.30 1.25 11.00 ;
        RECT  6.50 9.05 7.20 11.00 ;
        RECT  9.30 9.05 10.00 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.10 ;
        RECT  3.15 2.00 3.85 3.10 ;
        RECT  7.45 2.00 8.15 4.35 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 2.45 2.55 3.15 ;
        RECT  2.05 2.45 2.55 4.25 ;
        RECT  3.90 8.05 4.60 10.45 ;
        RECT  4.50 2.45 4.80 5.60 ;
        RECT  4.10 3.75 4.80 5.60 ;
        RECT  4.50 2.45 5.00 4.25 ;
        RECT  2.05 3.75 5.00 4.25 ;
        RECT  4.50 2.45 5.20 3.15 ;
        RECT  5.80 2.45 6.30 5.55 ;
        RECT  5.45 4.85 6.30 5.55 ;
        RECT  5.80 2.45 6.55 3.15 ;
        RECT  5.45 5.05 8.60 5.55 ;
        RECT  7.20 5.05 7.70 8.55 ;
        RECT  3.90 8.05 7.70 8.55 ;
        RECT  7.20 5.05 8.60 5.75 ;
    END
END OA32X2
MACRO OA32X4
    CLASS CORE ;
    FOREIGN OA32X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  8.15 6.70 8.65 10.55 ;
        RECT  7.95 8.95 8.65 10.55 ;
        RECT  8.70 2.75 9.40 4.35 ;
        RECT  8.90 2.75 9.40 7.60 ;
        RECT  8.15 6.70 9.55 7.60 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.35 7.60 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 6.70 6.75 7.60 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 4.00 7.60 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.60 8.20 1.30 11.00 ;
        RECT  6.60 9.00 7.30 11.00 ;
        RECT  9.30 8.20 10.00 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.10 ;
        RECT  3.15 2.00 3.85 3.10 ;
        RECT  7.35 2.00 8.05 4.35 ;
        RECT  10.05 2.00 10.75 4.35 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 2.45 2.55 3.15 ;
        RECT  2.05 2.45 2.55 4.25 ;
        RECT  3.95 8.05 4.65 10.45 ;
        RECT  4.50 2.45 4.80 5.55 ;
        RECT  4.10 3.75 4.80 5.55 ;
        RECT  4.50 2.45 5.00 4.25 ;
        RECT  2.05 3.75 5.00 4.25 ;
        RECT  4.50 2.45 5.20 3.15 ;
        RECT  5.80 2.45 6.30 5.55 ;
        RECT  5.45 4.80 6.30 5.55 ;
        RECT  5.80 2.45 6.55 3.15 ;
        RECT  5.45 5.05 8.45 5.55 ;
        RECT  7.20 5.05 7.70 8.55 ;
        RECT  3.95 8.05 7.70 8.55 ;
        RECT  7.20 5.05 8.45 5.75 ;
    END
END OA32X4
MACRO OA331X1
    CLASS CORE ;
    FOREIGN OA331X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.25 8.95 10.95 10.55 ;
        RECT  11.05 3.30 12.15 4.00 ;
        RECT  11.45 6.70 11.95 9.50 ;
        RECT  11.65 3.30 11.95 9.50 ;
        RECT  10.25 8.95 11.95 9.50 ;
        RECT  11.65 3.30 12.15 7.60 ;
        RECT  11.45 6.70 12.35 7.60 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.40 9.80 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  7.25 6.70 8.15 7.60 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  5.80 6.35 6.75 7.60 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  4.40 6.70 5.35 7.60 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.80 9.15 4.50 11.00 ;
        RECT  8.90 9.00 9.60 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.00 ;
        RECT  3.15 2.00 3.85 2.90 ;
        RECT  11.05 2.00 11.75 2.65 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  9.80 4.45 10.75 4.95 ;
        RECT  0.45 8.05 1.15 10.55 ;
        RECT  1.80 2.55 2.50 3.90 ;
        RECT  1.80 3.40 5.00 3.90 ;
        RECT  4.50 2.55 5.00 5.90 ;
        RECT  4.50 2.55 5.25 3.25 ;
        RECT  6.05 2.55 6.15 4.95 ;
        RECT  5.45 3.75 6.15 4.95 ;
        RECT  6.05 2.55 6.80 4.25 ;
        RECT  6.80 4.75 7.50 5.90 ;
        RECT  4.50 5.40 7.50 5.90 ;
        RECT  7.20 8.05 7.90 10.55 ;
        RECT  7.60 2.45 8.30 3.15 ;
        RECT  5.45 3.75 9.10 4.25 ;
        RECT  8.40 3.75 9.10 4.95 ;
        RECT  9.20 7.10 9.70 8.55 ;
        RECT  0.45 8.05 9.70 8.55 ;
        RECT  7.60 2.65 10.30 3.15 ;
        RECT  10.25 2.65 10.30 7.60 ;
        RECT  9.80 2.65 10.30 4.95 ;
        RECT  10.25 4.45 10.75 7.60 ;
        RECT  9.20 7.10 10.75 7.60 ;
        RECT  10.25 5.30 11.05 6.05 ;
    END
END OA331X1
MACRO OA331X2
    CLASS CORE ;
    FOREIGN OA331X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.25 8.05 10.95 10.55 ;
        RECT  11.45 2.75 12.15 4.45 ;
        RECT  11.45 6.70 11.95 8.55 ;
        RECT  11.65 2.75 11.95 8.55 ;
        RECT  10.25 8.05 11.95 8.55 ;
        RECT  11.65 2.75 12.15 7.60 ;
        RECT  11.45 6.70 12.35 7.60 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.40 9.80 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  7.25 6.70 8.15 7.60 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  5.80 6.35 6.75 7.60 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  4.40 6.70 5.35 7.60 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.80 9.15 4.50 11.00 ;
        RECT  8.90 9.00 9.60 11.00 ;
        RECT  11.60 9.00 12.30 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.00 ;
        RECT  3.15 2.00 3.85 2.90 ;
        RECT  12.80 2.00 13.50 4.45 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 8.05 1.15 10.55 ;
        RECT  1.80 2.55 2.50 3.90 ;
        RECT  1.80 3.40 5.00 3.90 ;
        RECT  4.50 2.55 5.00 5.90 ;
        RECT  4.50 2.55 5.25 3.25 ;
        RECT  6.05 2.55 6.15 4.95 ;
        RECT  5.45 3.75 6.15 4.95 ;
        RECT  6.05 2.55 6.80 4.25 ;
        RECT  6.80 4.75 7.50 5.90 ;
        RECT  4.50 5.40 7.50 5.90 ;
        RECT  7.20 8.05 7.90 10.55 ;
        RECT  7.60 2.45 8.30 3.15 ;
        RECT  5.45 3.75 9.10 4.25 ;
        RECT  8.40 3.75 9.10 4.95 ;
        RECT  9.20 7.10 9.70 8.55 ;
        RECT  0.45 8.05 9.70 8.55 ;
        RECT  7.60 2.65 10.75 3.15 ;
        RECT  10.25 2.65 10.75 7.60 ;
        RECT  9.20 7.10 10.75 7.60 ;
        RECT  10.25 5.30 11.20 6.00 ;
    END
END OA331X2
MACRO OA331X4
    CLASS CORE ;
    FOREIGN OA331X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.20 8.05 10.90 10.55 ;
        RECT  11.45 2.45 12.15 4.45 ;
        RECT  11.45 6.70 11.95 8.55 ;
        RECT  11.65 2.45 11.95 8.55 ;
        RECT  10.20 8.05 11.95 8.55 ;
        RECT  11.65 2.45 12.15 7.60 ;
        RECT  11.45 6.70 12.35 7.60 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.88 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.40 9.80 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  7.25 6.35 8.15 7.60 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  5.80 6.35 6.75 7.60 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  4.40 6.70 5.35 7.60 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.80 9.15 4.50 11.00 ;
        RECT  8.85 9.00 9.55 11.00 ;
        RECT  11.55 9.00 12.25 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.00 ;
        RECT  3.15 2.00 3.85 2.90 ;
        RECT  12.80 2.00 13.50 4.45 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 8.05 1.15 10.55 ;
        RECT  1.80 2.55 2.50 3.90 ;
        RECT  1.80 3.40 5.00 3.90 ;
        RECT  4.50 2.55 5.00 5.90 ;
        RECT  4.50 2.55 5.25 3.25 ;
        RECT  6.05 2.55 6.15 4.95 ;
        RECT  5.45 3.75 6.15 4.95 ;
        RECT  6.05 2.55 6.80 4.25 ;
        RECT  6.90 4.75 7.60 5.90 ;
        RECT  4.50 5.40 7.60 5.90 ;
        RECT  7.20 8.05 7.90 10.55 ;
        RECT  7.60 2.45 8.30 3.15 ;
        RECT  5.45 3.75 9.10 4.25 ;
        RECT  8.40 3.75 9.10 4.95 ;
        RECT  8.95 6.75 9.45 8.55 ;
        RECT  0.45 8.05 9.45 8.55 ;
        RECT  7.60 2.65 10.75 3.15 ;
        RECT  10.25 2.65 10.75 7.25 ;
        RECT  8.95 6.75 10.75 7.25 ;
        RECT  10.25 5.30 11.20 6.00 ;
    END
END OA331X4
MACRO OA332X1
    CLASS CORE ;
    FOREIGN OA332X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.20 8.85 11.90 10.45 ;
        RECT  12.85 2.45 13.35 9.35 ;
        RECT  11.20 8.85 13.35 9.35 ;
        RECT  12.85 2.45 13.55 3.15 ;
        RECT  12.85 6.70 13.75 7.60 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  8.65 6.70 9.55 7.60 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  7.25 6.70 8.15 7.60 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  5.85 6.35 6.75 7.60 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  4.10 9.40 4.80 11.00 ;
        RECT  9.80 9.00 10.50 11.00 ;
        RECT  12.85 10.05 13.55 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.00 ;
        RECT  3.15 2.00 3.85 2.70 ;
        RECT  11.50 2.00 12.20 3.15 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.70 4.20 7.85 4.30 ;
        RECT  0.75 8.05 1.45 10.00 ;
        RECT  1.80 2.55 2.50 3.70 ;
        RECT  4.50 2.55 5.20 3.70 ;
        RECT  1.80 3.20 5.20 3.70 ;
        RECT  4.70 2.55 5.20 4.30 ;
        RECT  0.75 8.05 5.90 8.55 ;
        RECT  5.40 8.05 5.90 9.35 ;
        RECT  5.80 4.75 6.50 5.85 ;
        RECT  5.85 2.60 6.55 3.30 ;
        RECT  7.15 3.80 7.65 4.90 ;
        RECT  4.70 3.80 7.65 4.30 ;
        RECT  7.15 4.20 7.85 4.90 ;
        RECT  5.85 2.60 8.80 3.10 ;
        RECT  7.45 8.85 8.15 10.45 ;
        RECT  7.95 2.60 8.80 3.30 ;
        RECT  8.25 8.05 8.75 9.35 ;
        RECT  5.40 8.85 8.75 9.35 ;
        RECT  8.30 2.60 8.80 5.85 ;
        RECT  5.80 5.35 8.80 5.85 ;
        RECT  8.30 4.35 9.30 5.05 ;
        RECT  9.30 2.60 10.60 3.30 ;
        RECT  10.10 2.60 10.60 8.55 ;
        RECT  8.25 8.05 10.60 8.55 ;
        RECT  10.10 4.80 10.80 5.50 ;
        RECT  10.10 7.60 11.85 8.30 ;
        RECT  8.25 8.05 11.85 8.30 ;
    END
END OA332X1
MACRO OA332X2
    CLASS CORE ;
    FOREIGN OA332X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.20 8.20 11.90 10.55 ;
        RECT  12.85 2.45 13.35 8.70 ;
        RECT  11.20 8.20 13.35 8.70 ;
        RECT  12.85 2.45 13.55 4.05 ;
        RECT  12.85 6.70 13.75 7.60 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  8.65 6.70 9.55 7.60 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  7.25 6.70 8.15 7.60 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  5.85 6.35 6.75 7.60 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  4.10 9.00 4.80 11.00 ;
        RECT  9.80 9.15 10.50 11.00 ;
        RECT  12.55 9.15 13.25 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.00 ;
        RECT  3.15 2.00 3.85 2.70 ;
        RECT  11.50 2.00 12.20 3.85 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.70 4.20 7.85 4.30 ;
        RECT  0.75 8.05 1.45 10.00 ;
        RECT  1.80 2.55 2.50 3.70 ;
        RECT  4.50 2.55 5.20 3.70 ;
        RECT  1.80 3.20 5.20 3.70 ;
        RECT  4.70 2.55 5.20 4.30 ;
        RECT  5.80 4.75 6.50 5.85 ;
        RECT  5.85 2.60 6.55 3.30 ;
        RECT  7.15 3.80 7.65 4.90 ;
        RECT  4.70 3.80 7.65 4.30 ;
        RECT  7.15 4.20 7.85 4.90 ;
        RECT  5.85 2.60 8.80 3.10 ;
        RECT  7.45 8.05 8.15 10.55 ;
        RECT  7.95 2.60 8.80 3.30 ;
        RECT  8.30 2.60 8.80 5.85 ;
        RECT  5.80 5.35 8.80 5.85 ;
        RECT  8.30 4.35 9.30 5.05 ;
        RECT  9.30 2.60 10.60 3.30 ;
        RECT  10.10 2.60 10.60 8.55 ;
        RECT  0.75 8.05 10.60 8.55 ;
        RECT  10.10 4.80 10.80 5.50 ;
        RECT  10.10 7.05 12.35 7.75 ;
    END
END OA332X2
MACRO OA332X4
    CLASS CORE ;
    FOREIGN OA332X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  11.50 8.20 12.20 10.55 ;
        RECT  12.85 2.45 13.35 8.70 ;
        RECT  11.50 8.20 13.35 8.70 ;
        RECT  12.70 2.45 13.40 4.35 ;
        RECT  12.85 6.70 13.75 7.60 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  8.65 6.50 9.55 7.60 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.23 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.35 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  7.25 6.70 8.15 7.60 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  5.85 6.35 6.75 7.60 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.35 7.60 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  0.25 6.70 1.15 7.60 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  4.30 9.00 5.00 11.00 ;
        RECT  10.15 9.15 10.85 11.00 ;
        RECT  12.85 9.15 13.55 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.00 ;
        RECT  3.15 2.00 3.85 2.70 ;
        RECT  11.35 2.00 12.05 3.85 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.70 4.20 7.65 4.30 ;
        RECT  9.90 4.80 10.60 5.50 ;
        RECT  0.85 8.05 1.55 10.00 ;
        RECT  1.80 2.55 2.50 3.70 ;
        RECT  4.50 2.55 5.20 3.70 ;
        RECT  1.80 3.20 5.20 3.70 ;
        RECT  4.70 2.55 5.20 4.30 ;
        RECT  5.60 4.75 6.30 5.85 ;
        RECT  5.85 2.60 6.55 3.30 ;
        RECT  6.95 3.80 7.45 4.90 ;
        RECT  4.70 3.80 7.45 4.30 ;
        RECT  6.95 4.20 7.65 4.90 ;
        RECT  5.85 2.60 8.60 3.10 ;
        RECT  7.75 2.60 8.60 3.30 ;
        RECT  7.65 8.05 8.35 10.05 ;
        RECT  8.10 2.60 8.60 5.85 ;
        RECT  5.60 5.35 8.60 5.85 ;
        RECT  8.10 4.35 9.10 5.05 ;
        RECT  9.10 2.60 10.40 3.30 ;
        RECT  10.10 2.60 10.40 8.55 ;
        RECT  9.90 2.60 10.40 5.50 ;
        RECT  10.10 4.80 10.60 8.55 ;
        RECT  0.85 8.05 10.60 8.55 ;
        RECT  11.70 7.05 12.40 7.75 ;
        RECT  10.10 7.25 12.40 7.75 ;
    END
END OA332X4
MACRO OA333X1
    CLASS CORE ;
    FOREIGN OA333X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  12.75 8.95 13.45 10.55 ;
        RECT  14.25 3.80 14.75 9.45 ;
        RECT  12.75 8.95 14.75 9.45 ;
        RECT  14.25 3.80 14.95 4.50 ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END Q
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  8.65 6.70 9.55 7.60 ;
        END
    END J
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  10.05 6.70 10.95 7.60 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  12.85 6.70 13.75 7.60 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 6.70 8.15 7.60 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 6.70 6.75 7.60 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.35 7.60 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.00 5.35 3.95 6.35 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.80 9.00 5.40 11.00 ;
        RECT  11.40 9.00 12.10 11.00 ;
        RECT  14.25 9.95 14.95 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.15 ;
        RECT  3.15 2.00 3.85 3.15 ;
        RECT  12.90 2.00 13.60 4.50 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 8.05 1.15 10.55 ;
        RECT  1.80 2.45 2.50 4.25 ;
        RECT  4.50 2.45 5.20 4.25 ;
        RECT  5.40 4.70 6.10 5.40 ;
        RECT  5.60 4.70 6.10 6.25 ;
        RECT  5.85 2.45 6.55 3.15 ;
        RECT  1.80 3.75 7.25 4.25 ;
        RECT  6.75 3.75 7.25 5.30 ;
        RECT  6.75 4.60 7.45 5.30 ;
        RECT  8.10 2.45 8.80 3.15 ;
        RECT  5.85 2.65 8.80 3.15 ;
        RECT  8.05 8.05 8.75 10.55 ;
        RECT  8.30 2.45 8.80 6.25 ;
        RECT  8.10 4.60 8.80 6.25 ;
        RECT  9.45 2.45 10.15 3.15 ;
        RECT  9.65 2.45 10.15 5.30 ;
        RECT  9.45 4.60 10.15 5.30 ;
        RECT  10.80 4.60 11.30 6.25 ;
        RECT  5.60 5.75 11.30 6.25 ;
        RECT  10.80 4.60 11.50 5.30 ;
        RECT  9.65 3.65 12.45 4.15 ;
        RECT  11.90 5.75 12.40 8.55 ;
        RECT  11.95 3.65 12.40 8.55 ;
        RECT  0.45 8.05 12.40 8.55 ;
        RECT  11.95 3.65 12.45 6.25 ;
        RECT  11.95 5.55 13.80 6.25 ;
        RECT  11.90 5.75 13.80 6.25 ;
    END
END OA333X1
MACRO OA333X2
    CLASS CORE ;
    FOREIGN OA333X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  12.75 8.05 13.45 10.55 ;
        RECT  14.25 2.80 14.75 8.55 ;
        RECT  12.75 8.05 14.75 8.55 ;
        RECT  14.25 2.80 14.95 4.50 ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END Q
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  8.65 6.70 9.55 7.60 ;
        END
    END J
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  10.05 6.70 10.95 7.60 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  12.85 6.70 13.75 7.60 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 6.70 8.15 7.60 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 6.70 6.75 7.60 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.35 7.60 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.00 5.35 3.95 6.35 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.80 9.00 5.40 11.00 ;
        RECT  11.40 9.00 12.10 11.00 ;
        RECT  14.10 9.00 14.80 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.15 ;
        RECT  3.15 2.00 3.85 3.15 ;
        RECT  12.90 2.00 13.60 4.50 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 8.05 1.15 10.55 ;
        RECT  1.80 2.45 2.50 4.25 ;
        RECT  4.50 2.45 5.20 4.25 ;
        RECT  5.40 4.70 6.10 5.40 ;
        RECT  5.60 4.70 6.10 6.25 ;
        RECT  5.85 2.45 6.55 3.15 ;
        RECT  1.80 3.75 7.25 4.25 ;
        RECT  6.75 3.75 7.25 5.30 ;
        RECT  6.75 4.60 7.45 5.30 ;
        RECT  8.10 2.45 8.80 3.15 ;
        RECT  5.85 2.65 8.80 3.15 ;
        RECT  8.05 8.05 8.75 10.55 ;
        RECT  8.30 2.45 8.80 6.25 ;
        RECT  8.10 4.60 8.80 6.25 ;
        RECT  9.45 2.45 10.15 3.15 ;
        RECT  9.65 2.45 10.15 5.30 ;
        RECT  9.45 4.60 10.15 5.30 ;
        RECT  10.80 4.60 11.30 6.25 ;
        RECT  5.60 5.75 11.30 6.25 ;
        RECT  10.80 4.60 11.50 5.30 ;
        RECT  9.65 3.65 12.45 4.15 ;
        RECT  11.80 5.75 12.30 8.55 ;
        RECT  11.95 3.65 12.30 8.55 ;
        RECT  0.45 8.05 12.30 8.55 ;
        RECT  11.95 3.65 12.45 6.25 ;
        RECT  11.95 5.55 13.80 6.25 ;
        RECT  11.80 5.75 13.80 6.25 ;
    END
END OA333X2
MACRO OA333X4
    CLASS CORE ;
    FOREIGN OA333X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  12.90 8.05 13.60 10.55 ;
        RECT  14.10 2.45 14.80 4.40 ;
        RECT  14.25 2.45 14.75 8.55 ;
        RECT  12.90 8.05 14.75 8.55 ;
        RECT  14.25 2.45 14.80 6.30 ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END Q
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  8.65 6.70 9.55 7.60 ;
        END
    END J
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  10.05 6.70 10.95 7.60 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  12.85 6.50 13.75 7.60 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 6.70 8.15 7.60 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 6.70 6.75 7.60 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.35 7.60 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.00 5.35 3.95 6.35 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.80 9.00 5.40 11.00 ;
        RECT  11.55 9.00 12.25 11.00 ;
        RECT  14.25 9.00 14.95 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.15 ;
        RECT  3.15 2.00 3.85 3.15 ;
        RECT  11.10 2.00 11.80 3.05 ;
        RECT  12.75 2.00 13.45 3.40 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 8.05 1.15 10.55 ;
        RECT  1.80 2.45 2.50 4.25 ;
        RECT  4.50 2.45 5.20 4.25 ;
        RECT  5.40 4.70 6.10 5.40 ;
        RECT  5.60 4.70 6.10 6.25 ;
        RECT  5.85 2.45 6.55 3.15 ;
        RECT  1.80 3.75 7.25 4.25 ;
        RECT  6.75 3.75 7.25 5.30 ;
        RECT  6.75 4.60 7.45 5.30 ;
        RECT  8.10 2.45 8.80 3.15 ;
        RECT  5.85 2.65 8.80 3.15 ;
        RECT  8.05 8.05 8.75 10.55 ;
        RECT  8.30 2.45 8.80 6.25 ;
        RECT  8.10 4.60 8.80 6.25 ;
        RECT  9.45 2.45 10.15 3.15 ;
        RECT  9.65 2.45 10.15 5.30 ;
        RECT  9.45 4.60 10.15 5.30 ;
        RECT  10.80 4.70 11.30 6.25 ;
        RECT  5.60 5.75 11.30 6.25 ;
        RECT  10.80 4.70 11.50 5.40 ;
        RECT  9.65 3.75 12.45 4.25 ;
        RECT  11.90 5.70 12.40 8.55 ;
        RECT  11.95 3.75 12.40 8.55 ;
        RECT  0.45 8.05 12.40 8.55 ;
        RECT  11.95 3.75 12.45 6.15 ;
        RECT  11.90 5.70 12.45 6.15 ;
        RECT  11.95 4.85 13.80 5.55 ;
    END
END OA333X4
MACRO OA33X1
    CLASS CORE ;
    FOREIGN OA33X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  9.45 4.10 10.95 4.40 ;
        RECT  10.25 3.70 10.50 10.55 ;
        RECT  9.45 3.70 10.50 4.40 ;
        RECT  10.25 4.10 10.75 10.55 ;
        RECT  10.05 8.95 10.75 10.55 ;
        RECT  10.05 4.10 10.95 5.00 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.35 7.60 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  7.00 6.70 8.15 7.60 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  8.65 6.70 9.55 7.60 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 8.40 1.15 11.00 ;
        RECT  8.70 9.10 9.40 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.05 ;
        RECT  3.15 2.00 3.85 3.05 ;
        RECT  9.45 2.00 10.15 2.95 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 3.65 7.85 4.10 ;
        RECT  1.80 2.45 2.55 4.10 ;
        RECT  3.80 8.10 4.50 9.70 ;
        RECT  4.50 2.45 5.15 5.35 ;
        RECT  4.45 3.60 5.15 5.35 ;
        RECT  4.50 2.45 5.20 4.15 ;
        RECT  1.80 3.60 5.20 4.10 ;
        RECT  5.10 8.10 5.80 9.70 ;
        RECT  5.80 4.60 6.30 8.60 ;
        RECT  3.80 8.10 6.30 8.60 ;
        RECT  5.80 4.60 6.50 6.25 ;
        RECT  5.85 2.45 6.55 3.20 ;
        RECT  4.45 3.65 7.85 4.15 ;
        RECT  7.15 3.65 7.85 5.30 ;
        RECT  5.85 2.70 9.00 3.20 ;
        RECT  8.30 2.70 8.80 6.25 ;
        RECT  5.80 5.75 8.80 6.25 ;
        RECT  8.30 2.70 9.00 3.45 ;
    END
END OA33X1
MACRO OA33X2
    CLASS CORE ;
    FOREIGN OA33X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.00 6.70 10.50 10.25 ;
        RECT  10.00 8.65 10.70 10.25 ;
        RECT  10.75 2.75 11.25 7.60 ;
        RECT  10.00 6.70 11.25 7.60 ;
        RECT  10.75 2.75 11.45 4.35 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.35 7.60 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  6.80 6.70 8.15 7.60 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  8.60 6.70 9.55 7.60 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 8.40 1.15 11.00 ;
        RECT  8.50 8.20 9.20 11.00 ;
        RECT  11.35 8.65 12.05 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.05 ;
        RECT  3.15 2.00 3.85 3.05 ;
        RECT  9.40 2.00 10.10 4.35 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 3.65 7.95 4.10 ;
        RECT  1.80 2.45 2.55 4.10 ;
        RECT  3.80 8.95 4.50 10.55 ;
        RECT  4.50 2.45 5.20 4.10 ;
        RECT  4.55 2.45 5.20 5.35 ;
        RECT  1.80 3.60 5.20 4.10 ;
        RECT  4.55 3.65 5.25 5.35 ;
        RECT  5.10 8.95 5.80 10.55 ;
        RECT  5.80 5.75 6.30 9.45 ;
        RECT  5.90 4.60 6.30 9.45 ;
        RECT  3.80 8.95 6.30 9.45 ;
        RECT  5.85 2.45 6.55 3.20 ;
        RECT  5.90 4.60 6.60 6.25 ;
        RECT  4.55 3.65 7.95 4.15 ;
        RECT  7.25 3.65 7.95 5.30 ;
        RECT  5.85 2.70 8.95 3.20 ;
        RECT  8.45 2.70 8.95 6.25 ;
        RECT  8.45 5.50 10.30 6.25 ;
        RECT  5.80 5.75 10.30 6.25 ;
    END
END OA33X2
MACRO OA33X4
    CLASS CORE ;
    FOREIGN OA33X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.50 2.75 11.20 4.35 ;
        RECT  10.25 6.70 10.75 10.55 ;
        RECT  10.70 2.75 10.75 10.55 ;
        RECT  10.05 8.05 10.75 10.55 ;
        RECT  10.05 9.30 10.95 10.20 ;
        RECT  10.70 2.75 11.20 7.20 ;
        RECT  10.25 6.70 11.20 7.20 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.35 7.60 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  6.85 6.70 7.75 7.40 ;
        RECT  7.25 6.70 7.75 8.90 ;
        RECT  7.25 8.00 8.15 8.90 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  8.30 6.70 9.55 7.45 ;
        RECT  8.65 6.70 9.55 7.60 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 8.05 1.15 11.00 ;
        RECT  8.70 8.05 9.40 11.00 ;
        RECT  11.40 8.05 12.10 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.05 ;
        RECT  3.15 2.00 3.85 3.05 ;
        RECT  9.15 2.00 9.85 4.35 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 2.45 2.50 4.15 ;
        RECT  3.80 8.95 4.50 10.55 ;
        RECT  4.50 2.45 5.00 5.30 ;
        RECT  4.30 3.65 5.00 5.30 ;
        RECT  4.50 2.45 5.20 4.15 ;
        RECT  5.65 4.60 6.35 5.30 ;
        RECT  5.80 4.60 5.85 10.55 ;
        RECT  5.15 8.95 5.85 10.55 ;
        RECT  5.80 4.60 6.30 9.45 ;
        RECT  3.80 8.95 6.30 9.45 ;
        RECT  5.80 4.60 6.35 6.25 ;
        RECT  5.85 2.45 6.55 3.20 ;
        RECT  1.80 3.65 7.70 4.15 ;
        RECT  7.00 3.65 7.70 5.30 ;
        RECT  5.85 2.70 8.65 3.20 ;
        RECT  8.15 2.70 8.65 6.25 ;
        RECT  9.55 5.50 10.25 6.25 ;
        RECT  5.80 5.75 10.25 6.25 ;
    END
END OA33X4
MACRO ON211X1
    CLASS CORE ;
    FOREIGN ON211X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.80 3.40 2.55 4.10 ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  2.00 3.40 2.55 7.65 ;
        RECT  2.00 7.15 3.50 7.65 ;
        RECT  2.80 7.15 3.50 10.55 ;
        RECT  2.80 8.05 6.15 8.55 ;
        RECT  5.65 8.05 6.15 10.55 ;
        RECT  5.65 8.95 6.35 10.55 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.35 7.60 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.00 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.45 1.15 11.00 ;
        RECT  4.30 9.00 5.00 11.00 ;
        RECT  7.20 9.60 7.90 11.00 ;
        RECT  0.00 11.00 8.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  5.50 2.00 6.20 4.45 ;
        RECT  7.15 2.00 7.85 4.50 ;
        RECT  0.00 0.00 8.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 2.45 1.15 4.05 ;
        RECT  0.45 2.45 3.85 2.95 ;
        RECT  3.15 2.45 3.85 4.05 ;
    END
END ON211X1
MACRO ON211X2
    CLASS CORE ;
    FOREIGN ON211X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.80 3.40 2.50 4.10 ;
        RECT  4.50 3.40 5.35 4.10 ;
        RECT  1.80 3.60 5.35 4.10 ;
        RECT  4.45 5.40 5.35 6.30 ;
        RECT  4.80 3.40 5.35 7.75 ;
        RECT  4.80 7.05 8.05 7.75 ;
        RECT  7.35 7.05 8.05 10.55 ;
        RECT  4.80 7.05 10.75 7.60 ;
        RECT  10.05 7.05 10.75 10.55 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.50 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 11.00 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.50 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.25 9.55 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.88 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.88 ;
        PORT
        LAYER M1M ;
        RECT  5.80 5.40 6.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 9.55 2.45 11.00 ;
        RECT  3.25 7.10 3.95 11.00 ;
        RECT  3.25 9.40 5.70 10.10 ;
        RECT  8.70 8.05 9.40 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  10.75 2.00 11.45 4.45 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 2.45 1.15 4.25 ;
        RECT  3.15 2.45 3.85 3.15 ;
        RECT  0.45 2.45 6.55 2.95 ;
        RECT  5.85 2.45 6.55 4.45 ;
        RECT  5.85 3.75 9.10 4.45 ;
    END
END ON211X2
MACRO ON211X4
    CLASS CORE ;
    FOREIGN ON211X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.80 3.40 2.50 4.10 ;
        RECT  4.50 3.40 5.20 4.10 ;
        RECT  7.20 3.40 7.90 4.10 ;
        RECT  5.20 9.15 11.65 9.85 ;
        RECT  9.90 3.40 10.60 4.10 ;
        RECT  1.80 3.60 10.60 4.10 ;
        RECT  10.10 3.40 10.60 7.60 ;
        RECT  10.05 9.15 11.65 10.20 ;
        RECT  10.95 7.10 11.65 10.55 ;
        RECT  18.60 7.10 19.30 10.55 ;
        RECT  10.10 7.10 22.00 7.60 ;
        RECT  21.30 7.10 22.00 10.55 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 7.00 ;
        PORT
        LAYER M1M ;
        RECT  21.25 5.40 22.40 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 7.00 ;
        PORT
        LAYER M1M ;
        RECT  19.50 5.40 20.75 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.40 9.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  11.05 5.40 12.35 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 9.60 2.05 11.00 ;
        RECT  2.85 7.00 3.55 11.00 ;
        RECT  4.45 6.80 7.95 7.50 ;
        RECT  2.85 7.00 7.95 7.50 ;
        RECT  12.60 8.05 16.00 11.00 ;
        RECT  17.25 8.05 17.95 11.00 ;
        RECT  19.95 8.05 20.65 11.00 ;
        RECT  22.65 8.05 23.35 11.00 ;
        RECT  0.00 11.00 23.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  22.15 2.00 22.85 4.45 ;
        RECT  0.00 0.00 23.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 2.45 1.15 4.10 ;
        RECT  3.15 2.45 3.85 3.15 ;
        RECT  5.85 2.45 6.55 3.15 ;
        RECT  8.55 2.45 9.25 3.15 ;
        RECT  0.45 2.45 11.95 2.95 ;
        RECT  11.25 2.45 11.95 4.25 ;
        RECT  11.25 3.55 20.50 4.25 ;
    END
END ON211X4
MACRO ON21X1
    CLASS CORE ;
    FOREIGN ON21X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.45 2.55 4.15 ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  2.05 2.45 2.55 7.80 ;
        RECT  2.05 7.25 4.20 7.80 ;
        RECT  3.50 7.25 4.20 10.25 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 9.55 1.15 11.00 ;
        RECT  2.00 9.40 2.70 11.00 ;
        RECT  5.85 7.25 6.55 11.00 ;
        RECT  0.00 11.00 7.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  4.50 2.00 5.20 4.00 ;
        RECT  0.00 0.00 7.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.15 2.45 3.85 4.95 ;
        RECT  5.85 2.45 6.55 4.95 ;
        RECT  3.15 4.45 6.55 4.95 ;
    END
END ON21X1
MACRO ON21X2
    CLASS CORE ;
    FOREIGN ON21X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.60 2.80 1.15 6.30 ;
        RECT  0.25 5.40 1.15 6.30 ;
        RECT  0.65 2.80 1.15 7.80 ;
        RECT  0.60 2.80 1.30 4.50 ;
        RECT  0.65 7.25 3.30 7.80 ;
        RECT  2.60 7.25 3.30 10.55 ;
        RECT  2.60 9.20 5.10 9.90 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.80 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.20 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.20 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.25 8.50 1.95 11.00 ;
        RECT  6.75 7.25 7.45 11.00 ;
        RECT  0.00 11.00 8.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.30 2.00 4.00 3.95 ;
        RECT  6.35 2.00 7.95 4.50 ;
        RECT  0.00 0.00 8.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.95 2.45 2.65 4.90 ;
        RECT  4.65 2.45 5.35 4.90 ;
        RECT  1.95 4.40 5.35 4.90 ;
    END
END ON21X2
MACRO ON21X4
    CLASS CORE ;
    FOREIGN ON21X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  2.05 3.40 2.50 10.55 ;
        RECT  1.80 3.40 2.50 6.30 ;
        RECT  2.05 4.60 2.55 10.55 ;
        RECT  2.05 8.05 2.75 10.55 ;
        RECT  2.05 8.05 5.45 8.60 ;
        RECT  4.50 3.40 5.20 5.10 ;
        RECT  1.80 4.60 5.20 5.10 ;
        RECT  4.75 8.05 5.45 10.55 ;
        RECT  4.75 9.15 11.10 9.85 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.60 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 8.40 ;
        PORT
        LAYER M1M ;
        RECT  11.10 5.40 12.35 6.35 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 8.40 ;
        PORT
        LAYER M1M ;
        RECT  5.05 5.75 5.55 7.60 ;
        RECT  4.45 6.70 5.55 7.60 ;
        RECT  5.05 5.75 5.90 6.45 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 9.55 1.15 11.00 ;
        RECT  3.40 9.05 4.10 11.00 ;
        RECT  7.10 6.80 13.45 7.50 ;
        RECT  12.75 6.80 13.45 11.00 ;
        RECT  14.25 9.55 14.95 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  7.50 2.00 8.20 3.95 ;
        RECT  10.20 2.00 10.90 3.95 ;
        RECT  12.90 2.00 13.60 3.95 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 2.45 1.15 4.15 ;
        RECT  3.15 2.45 3.85 4.15 ;
        RECT  0.45 2.45 6.85 2.95 ;
        RECT  6.15 2.45 6.85 4.90 ;
        RECT  8.85 2.45 9.55 4.90 ;
        RECT  11.55 2.45 12.25 4.90 ;
        RECT  14.25 2.45 14.95 4.90 ;
        RECT  6.15 4.40 14.95 4.90 ;
    END
END ON21X4
MACRO ON221X1
    CLASS CORE ;
    FOREIGN ON221X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.95 7.50 1.65 10.00 ;
        RECT  5.65 7.50 6.35 10.10 ;
        RECT  7.20 2.85 7.75 8.00 ;
        RECT  0.95 7.50 7.75 8.00 ;
        RECT  7.20 2.85 7.90 5.00 ;
        RECT  7.20 4.10 8.15 5.00 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.40 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.35 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.00 5.40 3.95 6.35 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.30 8.45 4.00 11.00 ;
        RECT  7.15 8.45 7.85 11.00 ;
        RECT  8.65 9.55 9.35 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.15 2.00 3.85 2.70 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 2.45 1.15 4.60 ;
        RECT  1.80 2.95 2.50 3.65 ;
        RECT  4.50 2.95 5.20 3.65 ;
        RECT  1.80 3.15 5.20 3.65 ;
        RECT  5.85 2.45 6.55 4.60 ;
        RECT  0.45 4.10 6.55 4.60 ;
    END
END ON221X1
MACRO ON221X2
    CLASS CORE ;
    FOREIGN ON221X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 18.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  2.30 6.90 3.00 9.60 ;
        RECT  11.90 6.90 12.60 9.60 ;
        RECT  14.80 6.90 15.50 10.55 ;
        RECT  15.65 5.40 16.15 7.40 ;
        RECT  2.30 6.90 16.15 7.40 ;
        RECT  15.65 5.40 16.55 6.30 ;
        RECT  14.15 2.45 17.40 3.15 ;
        RECT  16.70 2.45 17.20 5.90 ;
        RECT  15.65 5.40 17.20 5.90 ;
        RECT  16.70 2.45 17.40 4.50 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.50 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.20 6.40 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.30 12.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.30 2.55 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.35 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.35 6.75 6.35 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  5.00 8.80 5.70 11.00 ;
        RECT  9.20 8.80 9.90 11.00 ;
        RECT  16.15 7.85 16.85 11.00 ;
        RECT  0.00 11.00 18.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  4.60 2.00 5.30 2.40 ;
        RECT  7.30 2.00 8.00 2.40 ;
        RECT  0.00 0.00 18.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.55 2.45 1.25 4.05 ;
        RECT  0.95 7.70 1.65 10.55 ;
        RECT  1.90 3.40 2.60 4.60 ;
        RECT  3.25 2.45 3.95 3.35 ;
        RECT  0.55 2.45 3.95 2.95 ;
        RECT  3.65 7.85 4.35 10.55 ;
        RECT  0.95 10.05 4.35 10.55 ;
        RECT  3.65 7.85 7.05 8.35 ;
        RECT  5.95 2.65 6.65 3.35 ;
        RECT  6.35 7.85 7.05 10.55 ;
        RECT  7.85 7.85 8.55 10.55 ;
        RECT  8.65 2.45 9.35 3.35 ;
        RECT  3.25 2.85 9.35 3.35 ;
        RECT  7.85 7.85 11.25 8.35 ;
        RECT  10.00 3.40 10.70 4.60 ;
        RECT  10.55 7.85 11.25 10.55 ;
        RECT  8.65 2.45 12.05 2.95 ;
        RECT  0.55 2.85 12.05 2.95 ;
        RECT  11.35 2.45 12.05 3.15 ;
        RECT  12.85 2.45 13.55 4.60 ;
        RECT  13.25 7.85 13.95 10.55 ;
        RECT  10.55 10.05 13.95 10.55 ;
        RECT  12.85 3.80 16.05 4.60 ;
        RECT  1.90 4.10 16.05 4.60 ;
    END
END ON221X2
MACRO ON221X4
    CLASS CORE ;
    FOREIGN ON221X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 30.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  7.20 6.75 7.90 9.60 ;
        RECT  9.90 6.75 10.60 9.60 ;
        RECT  19.50 6.75 20.20 9.60 ;
        RECT  22.20 6.75 22.90 9.60 ;
        RECT  25.45 3.65 25.60 7.25 ;
        RECT  24.90 3.65 25.60 4.40 ;
        RECT  25.45 3.90 25.95 7.25 ;
        RECT  25.45 5.40 26.35 7.25 ;
        RECT  7.20 6.75 27.10 7.25 ;
        RECT  26.40 6.75 27.10 10.55 ;
        RECT  27.60 3.65 28.30 4.40 ;
        RECT  24.90 3.90 28.30 4.40 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 7.00 ;
        PORT
        LAYER M1M ;
        RECT  26.85 5.40 27.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.40 9.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.70 2.50 11.00 ;
        RECT  4.50 7.70 5.20 11.00 ;
        RECT  14.10 8.65 14.80 11.00 ;
        RECT  16.80 8.65 17.50 11.00 ;
        RECT  25.05 7.70 25.75 11.00 ;
        RECT  27.75 7.70 28.45 11.00 ;
        RECT  29.45 9.60 30.15 11.00 ;
        RECT  0.00 11.00 30.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 3.85 ;
        RECT  4.50 2.00 5.20 3.85 ;
        RECT  7.20 2.00 7.90 3.85 ;
        RECT  9.90 2.00 10.60 3.85 ;
        RECT  0.00 0.00 30.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 2.45 1.15 4.80 ;
        RECT  0.45 6.75 1.15 10.55 ;
        RECT  3.15 2.45 3.85 4.80 ;
        RECT  3.15 6.75 3.85 10.55 ;
        RECT  0.45 6.75 6.55 7.25 ;
        RECT  5.85 2.45 6.55 4.80 ;
        RECT  5.85 6.75 6.55 10.55 ;
        RECT  8.55 2.45 9.25 4.80 ;
        RECT  8.55 7.70 9.25 10.55 ;
        RECT  11.25 2.45 11.95 4.80 ;
        RECT  0.45 4.30 11.95 4.80 ;
        RECT  11.25 7.70 11.95 10.55 ;
        RECT  5.85 10.05 11.95 10.55 ;
        RECT  12.60 3.65 13.30 4.40 ;
        RECT  12.75 7.70 13.45 10.55 ;
        RECT  13.95 2.45 14.65 3.15 ;
        RECT  15.30 3.65 16.00 4.40 ;
        RECT  15.45 7.70 16.15 10.55 ;
        RECT  16.65 2.45 17.35 3.15 ;
        RECT  12.75 7.70 18.85 8.20 ;
        RECT  18.00 3.65 18.70 4.40 ;
        RECT  18.15 7.70 18.85 10.55 ;
        RECT  19.35 2.45 20.05 3.15 ;
        RECT  20.70 3.65 21.40 4.40 ;
        RECT  20.85 7.70 21.55 10.55 ;
        RECT  11.25 2.45 22.75 2.95 ;
        RECT  22.05 2.45 22.75 3.15 ;
        RECT  23.55 2.70 24.25 4.40 ;
        RECT  12.60 3.90 24.25 4.40 ;
        RECT  23.55 7.70 24.25 10.55 ;
        RECT  18.15 10.05 24.25 10.55 ;
        RECT  26.25 2.70 26.95 3.40 ;
        RECT  23.55 2.70 29.65 3.20 ;
        RECT  28.95 2.70 29.65 4.40 ;
    END
END ON221X4
MACRO ON222X1
    CLASS CORE ;
    FOREIGN ON222X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.95 8.05 7.70 8.35 ;
        RECT  0.95 7.85 1.65 10.55 ;
        RECT  4.55 7.85 5.05 8.55 ;
        RECT  0.95 7.85 5.05 8.35 ;
        RECT  5.65 8.05 6.35 10.55 ;
        RECT  7.20 3.55 7.70 8.55 ;
        RECT  4.55 8.05 7.70 8.55 ;
        RECT  7.20 3.55 7.90 4.25 ;
        RECT  7.20 5.40 8.15 6.30 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  8.65 6.70 9.55 7.60 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  5.85 6.70 6.75 7.60 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        RECT  4.45 5.40 5.65 6.20 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.35 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.35 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.30 8.80 4.00 11.00 ;
        RECT  8.00 9.00 8.70 11.00 ;
        RECT  9.80 9.55 10.50 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.15 2.00 3.85 3.05 ;
        RECT  10.05 2.00 10.75 4.70 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 2.55 1.15 4.95 ;
        RECT  1.80 3.30 2.50 4.00 ;
        RECT  4.50 3.30 5.20 4.00 ;
        RECT  1.80 3.50 5.20 4.00 ;
        RECT  5.85 2.55 6.55 4.95 ;
        RECT  0.45 4.45 6.55 4.95 ;
        RECT  5.85 2.55 9.25 3.05 ;
        RECT  8.55 2.55 9.25 4.35 ;
    END
END ON222X1
MACRO ON222X2
    CLASS CORE ;
    FOREIGN ON222X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  2.30 6.90 3.00 9.60 ;
        RECT  11.90 6.90 12.60 9.60 ;
        RECT  2.30 6.90 16.85 7.40 ;
        RECT  15.65 5.40 16.85 6.30 ;
        RECT  16.35 3.80 16.85 9.60 ;
        RECT  16.15 6.90 16.85 9.60 ;
        RECT  13.85 3.80 19.20 4.50 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.40 19.45 6.35 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.20 6.40 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.30 12.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.30 2.55 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.35 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.35 6.75 6.35 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  5.00 8.80 5.70 11.00 ;
        RECT  9.20 8.80 9.90 11.00 ;
        RECT  18.85 8.40 19.55 11.00 ;
        RECT  0.00 11.00 22.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  4.60 2.00 5.30 2.40 ;
        RECT  7.30 2.00 8.00 2.40 ;
        RECT  21.25 2.00 21.95 4.55 ;
        RECT  0.00 0.00 22.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.55 2.45 1.25 4.05 ;
        RECT  0.95 7.70 1.65 10.55 ;
        RECT  1.90 3.40 2.60 4.60 ;
        RECT  3.25 2.45 3.95 3.35 ;
        RECT  0.55 2.45 3.95 2.95 ;
        RECT  3.65 7.85 4.35 10.55 ;
        RECT  0.95 10.05 4.35 10.55 ;
        RECT  3.65 7.85 7.05 8.35 ;
        RECT  5.95 2.65 6.65 3.35 ;
        RECT  6.35 7.85 7.05 10.55 ;
        RECT  7.85 7.85 8.55 10.55 ;
        RECT  8.65 2.45 9.35 3.35 ;
        RECT  3.25 2.85 9.35 3.35 ;
        RECT  7.85 7.85 11.25 8.35 ;
        RECT  10.00 3.40 10.70 4.60 ;
        RECT  10.55 7.85 11.25 10.55 ;
        RECT  8.65 2.45 12.05 2.95 ;
        RECT  0.55 2.85 12.05 2.95 ;
        RECT  11.35 2.45 12.05 3.15 ;
        RECT  12.70 2.45 13.20 4.60 ;
        RECT  1.90 4.10 13.20 4.60 ;
        RECT  13.25 7.85 13.95 10.55 ;
        RECT  10.55 10.05 13.95 10.55 ;
        RECT  14.80 7.85 15.50 10.55 ;
        RECT  12.70 2.45 15.70 3.15 ;
        RECT  12.70 2.45 20.20 2.95 ;
        RECT  17.50 7.45 18.20 10.55 ;
        RECT  14.80 10.05 18.20 10.55 ;
        RECT  17.50 7.45 20.90 7.95 ;
        RECT  17.35 2.45 20.20 3.15 ;
        RECT  20.20 7.45 20.90 10.55 ;
    END
END ON222X2
MACRO ON222X4
    CLASS CORE ;
    FOREIGN ON222X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 37.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  7.20 6.75 7.90 9.60 ;
        RECT  9.90 6.75 10.60 9.60 ;
        RECT  19.50 6.75 20.20 9.60 ;
        RECT  22.20 6.75 22.90 9.60 ;
        RECT  24.90 3.65 25.60 4.40 ;
        RECT  27.60 3.65 28.30 4.40 ;
        RECT  29.65 3.90 30.15 7.25 ;
        RECT  29.65 5.40 30.55 7.25 ;
        RECT  30.30 3.65 31.00 4.40 ;
        RECT  31.80 6.75 32.50 9.60 ;
        RECT  33.00 3.65 33.70 4.40 ;
        RECT  24.90 3.90 33.70 4.40 ;
        RECT  7.20 6.75 35.20 7.25 ;
        RECT  34.50 6.75 35.20 9.60 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  26.85 5.40 27.75 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  32.45 5.40 33.35 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.40 9.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 7.70 2.50 11.00 ;
        RECT  4.50 7.70 5.20 11.00 ;
        RECT  14.10 8.65 14.80 11.00 ;
        RECT  16.80 8.65 17.50 11.00 ;
        RECT  26.40 8.65 27.10 11.00 ;
        RECT  29.10 8.65 29.80 11.00 ;
        RECT  0.00 11.00 37.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 3.85 ;
        RECT  4.50 2.00 5.20 3.85 ;
        RECT  7.20 2.00 7.90 3.85 ;
        RECT  9.90 2.00 10.60 3.85 ;
        RECT  36.25 2.00 36.95 4.40 ;
        RECT  0.00 0.00 37.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 2.45 1.15 4.80 ;
        RECT  0.45 6.75 1.15 10.55 ;
        RECT  3.15 2.45 3.85 4.80 ;
        RECT  3.15 6.75 3.85 10.55 ;
        RECT  0.45 6.75 6.55 7.25 ;
        RECT  5.85 2.45 6.55 4.80 ;
        RECT  5.85 6.75 6.55 10.55 ;
        RECT  8.55 2.45 9.25 4.80 ;
        RECT  8.55 7.70 9.25 10.55 ;
        RECT  11.25 2.45 11.95 4.80 ;
        RECT  0.45 4.30 11.95 4.80 ;
        RECT  11.25 7.70 11.95 10.55 ;
        RECT  5.85 10.05 11.95 10.55 ;
        RECT  12.60 3.65 13.30 4.40 ;
        RECT  12.75 7.70 13.45 10.55 ;
        RECT  13.95 2.45 14.65 3.15 ;
        RECT  15.30 3.65 16.00 4.40 ;
        RECT  15.45 7.70 16.15 10.55 ;
        RECT  16.65 2.45 17.35 3.15 ;
        RECT  12.75 7.70 18.85 8.20 ;
        RECT  18.00 3.65 18.70 4.40 ;
        RECT  18.15 7.70 18.85 10.55 ;
        RECT  19.35 2.45 20.05 3.15 ;
        RECT  20.70 3.65 21.40 4.40 ;
        RECT  20.85 7.70 21.55 10.55 ;
        RECT  11.25 2.45 22.75 2.95 ;
        RECT  22.05 2.45 22.75 3.15 ;
        RECT  23.55 2.70 24.25 4.40 ;
        RECT  12.60 3.90 24.25 4.40 ;
        RECT  23.55 7.70 24.25 10.55 ;
        RECT  18.15 10.05 24.25 10.55 ;
        RECT  25.05 7.70 25.75 10.55 ;
        RECT  26.25 2.70 26.95 3.40 ;
        RECT  27.75 7.70 28.45 10.55 ;
        RECT  28.95 2.70 29.65 3.40 ;
        RECT  25.05 7.70 31.15 8.20 ;
        RECT  30.45 7.70 31.15 10.55 ;
        RECT  31.65 2.70 32.35 3.40 ;
        RECT  33.15 7.70 33.85 10.55 ;
        RECT  23.55 2.70 35.05 3.20 ;
        RECT  34.35 2.70 35.05 4.40 ;
        RECT  35.85 7.70 36.55 10.55 ;
        RECT  30.45 10.05 36.55 10.55 ;
    END
END ON222X4
MACRO ON22X1
    CLASS CORE ;
    FOREIGN ON22X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  2.95 6.90 3.65 10.45 ;
        RECT  4.45 3.40 4.95 7.40 ;
        RECT  2.95 6.90 4.95 7.40 ;
        RECT  4.45 3.40 5.20 4.10 ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.35 2.55 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 8.15 1.15 11.00 ;
        RECT  5.30 7.85 6.00 11.00 ;
        RECT  0.00 11.00 7.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 3.20 ;
        RECT  0.00 0.00 7.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 2.45 1.15 4.15 ;
        RECT  3.10 2.45 3.85 4.15 ;
        RECT  0.45 3.65 3.85 4.15 ;
        RECT  3.10 2.45 6.55 2.95 ;
        RECT  5.85 2.45 6.55 4.10 ;
    END
END ON22X1
MACRO ON22X2
    CLASS CORE ;
    FOREIGN ON22X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.65 3.40 5.15 10.55 ;
        RECT  4.55 6.70 5.25 10.55 ;
        RECT  4.45 6.70 5.35 7.60 ;
        RECT  4.65 3.40 5.40 4.10 ;
        RECT  2.80 9.15 7.00 9.85 ;
        RECT  7.40 3.40 7.90 7.60 ;
        RECT  4.45 7.10 7.90 7.60 ;
        RECT  7.40 3.40 8.10 4.10 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.20 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.20 ;
        PORT
        LAYER M1M ;
        RECT  3.00 5.30 3.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.20 ;
        PORT
        LAYER M1M ;
        RECT  8.55 5.40 9.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.20 ;
        PORT
        LAYER M1M ;
        RECT  5.70 5.30 6.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.15 1.15 11.00 ;
        RECT  8.65 7.15 9.35 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.00 2.00 2.70 3.50 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.65 2.45 1.35 4.45 ;
        RECT  3.30 2.45 4.05 4.45 ;
        RECT  0.65 3.95 4.05 4.45 ;
        RECT  6.05 2.45 6.75 4.10 ;
        RECT  3.30 2.45 9.45 2.95 ;
        RECT  8.75 2.45 9.45 4.10 ;
    END
END ON22X2
MACRO ON22X4
    CLASS CORE ;
    FOREIGN ON22X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.35 4.80 10.85 10.55 ;
        RECT  10.65 3.65 10.85 10.55 ;
        RECT  10.15 6.85 10.85 10.55 ;
        RECT  10.05 9.15 10.95 10.55 ;
        RECT  10.65 3.65 11.15 5.30 ;
        RECT  10.35 4.80 11.15 5.30 ;
        RECT  13.10 3.40 13.80 4.15 ;
        RECT  15.80 3.40 16.50 4.15 ;
        RECT  4.50 9.15 16.50 9.85 ;
        RECT  18.50 3.40 19.20 4.15 ;
        RECT  10.65 3.65 19.20 4.15 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 8.40 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.35 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 8.40 ;
        PORT
        LAYER M1M ;
        RECT  7.65 4.80 8.15 6.30 ;
        RECT  7.25 5.40 8.15 6.30 ;
        RECT  7.65 4.80 8.35 5.50 ;
        RECT  7.25 5.40 8.35 5.50 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 8.40 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.35 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 8.40 ;
        PORT
        LAYER M1M ;
        RECT  12.65 5.40 13.75 5.50 ;
        RECT  12.85 4.80 13.40 6.30 ;
        RECT  12.65 4.80 13.40 5.50 ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.55 9.55 1.25 11.00 ;
        RECT  2.15 6.80 2.85 11.00 ;
        RECT  2.15 6.80 8.35 7.50 ;
        RECT  12.65 6.80 18.85 7.50 ;
        RECT  18.15 6.80 18.85 11.00 ;
        RECT  19.75 9.55 20.45 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.30 ;
        RECT  3.15 2.00 3.85 3.30 ;
        RECT  5.85 2.00 6.55 3.30 ;
        RECT  8.55 2.00 9.25 3.30 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 2.45 2.50 4.25 ;
        RECT  4.50 2.45 5.20 4.25 ;
        RECT  7.20 2.45 7.90 4.25 ;
        RECT  9.70 2.45 10.20 4.25 ;
        RECT  1.80 3.75 10.20 4.25 ;
        RECT  11.75 2.45 12.45 3.15 ;
        RECT  14.45 2.45 15.15 3.15 ;
        RECT  17.15 2.45 17.85 3.15 ;
        RECT  9.70 2.45 20.55 2.95 ;
        RECT  19.85 2.45 20.55 3.15 ;
    END
END ON22X4
MACRO ON311X1
    CLASS CORE ;
    FOREIGN ON311X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.20 6.30 ;
        RECT  0.70 5.40 1.20 8.80 ;
        RECT  1.50 8.30 2.20 10.05 ;
        RECT  2.25 2.85 2.75 5.90 ;
        RECT  0.25 5.40 2.75 5.90 ;
        RECT  2.25 2.85 2.95 4.45 ;
        RECT  0.70 8.30 6.00 8.80 ;
        RECT  4.20 8.30 4.90 10.05 ;
        RECT  5.30 7.15 6.00 8.85 ;
        RECT  4.20 8.30 6.00 8.85 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  1.65 6.70 2.55 7.60 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  3.05 6.70 3.95 7.60 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.70 6.35 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  6.95 5.25 8.15 5.95 ;
        RECT  7.25 5.25 8.15 6.35 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.40 9.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.85 9.40 3.55 11.00 ;
        RECT  8.65 7.15 9.35 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.60 2.00 1.30 4.50 ;
        RECT  5.95 2.00 6.65 3.40 ;
        RECT  8.65 2.00 9.35 4.45 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.60 2.55 5.30 4.45 ;
        RECT  7.30 2.55 8.00 4.45 ;
        RECT  4.60 3.95 8.00 4.45 ;
    END
END ON311X1
MACRO ON311X2
    CLASS CORE ;
    FOREIGN ON311X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        RECT  2.50 7.10 3.20 10.55 ;
        RECT  1.60 2.85 4.40 3.55 ;
        RECT  3.70 2.85 4.40 4.45 ;
        RECT  3.70 3.95 4.95 4.45 ;
        RECT  2.50 7.10 5.90 7.60 ;
        RECT  4.85 3.95 4.95 7.60 ;
        RECT  4.45 3.95 4.95 6.30 ;
        RECT  5.20 5.40 5.35 10.55 ;
        RECT  4.85 5.40 5.35 7.60 ;
        RECT  5.20 7.10 5.90 10.55 ;
        RECT  12.30 7.15 13.00 8.75 ;
        RECT  5.20 8.05 13.00 8.75 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.50 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 4.00 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.50 ;
        PORT
        LAYER M1M ;
        RECT  5.80 5.40 6.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  9.90 5.40 10.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.25 12.75 6.35 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 9.60 1.15 11.00 ;
        RECT  3.85 8.05 4.55 11.00 ;
        RECT  15.65 7.15 16.35 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 5.15 ;
        RECT  0.45 4.45 2.05 5.15 ;
        RECT  7.55 2.00 8.25 3.55 ;
        RECT  10.25 2.00 10.95 3.55 ;
        RECT  12.95 2.00 13.65 3.55 ;
        RECT  15.65 2.00 16.35 3.55 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  6.05 2.45 6.75 4.50 ;
        RECT  8.90 2.45 9.60 4.50 ;
        RECT  11.60 2.55 12.30 4.50 ;
        RECT  14.30 2.55 15.00 4.50 ;
        RECT  6.05 4.00 15.00 4.50 ;
    END
END ON311X2
MACRO ON311X4
    CLASS CORE ;
    FOREIGN ON311X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 30.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  16.95 6.75 17.65 9.60 ;
        RECT  19.65 6.75 20.35 9.60 ;
        RECT  22.35 6.75 23.05 10.55 ;
        RECT  25.45 3.40 25.65 10.55 ;
        RECT  24.95 3.40 25.65 4.10 ;
        RECT  25.45 3.60 25.75 10.55 ;
        RECT  25.05 6.75 25.75 10.55 ;
        RECT  25.45 3.60 25.95 7.25 ;
        RECT  25.45 5.40 26.35 7.25 ;
        RECT  16.95 6.75 28.45 7.25 ;
        RECT  27.65 3.40 28.35 4.10 ;
        RECT  24.95 3.60 28.35 4.10 ;
        RECT  27.75 6.75 28.45 10.55 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 7.00 ;
        PORT
        LAYER M1M ;
        RECT  26.85 5.40 27.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 7.00 ;
        PORT
        LAYER M1M ;
        RECT  22.65 5.40 23.55 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.65 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.55 9.55 1.25 11.00 ;
        RECT  2.10 7.15 2.80 11.00 ;
        RECT  4.80 7.70 5.50 11.00 ;
        RECT  7.50 7.70 8.20 11.00 ;
        RECT  23.70 7.70 24.40 11.00 ;
        RECT  26.40 7.70 27.10 11.00 ;
        RECT  29.45 9.60 30.15 11.00 ;
        RECT  0.00 11.00 30.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 3.60 ;
        RECT  4.50 2.00 5.20 3.60 ;
        RECT  7.20 2.00 7.90 3.60 ;
        RECT  9.90 2.00 10.60 3.60 ;
        RECT  12.60 2.00 13.30 3.60 ;
        RECT  15.30 2.00 16.00 3.60 ;
        RECT  0.00 0.00 30.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 2.45 1.15 4.60 ;
        RECT  3.15 2.45 3.85 4.60 ;
        RECT  3.45 6.75 4.15 10.55 ;
        RECT  5.85 2.45 6.55 4.60 ;
        RECT  6.15 6.75 6.85 10.55 ;
        RECT  3.45 6.75 9.55 7.25 ;
        RECT  8.55 2.45 9.25 4.60 ;
        RECT  8.85 6.75 9.55 10.55 ;
        RECT  10.20 6.75 10.90 9.60 ;
        RECT  11.25 2.45 11.95 4.60 ;
        RECT  11.55 7.70 12.25 10.55 ;
        RECT  12.90 6.75 13.60 9.60 ;
        RECT  13.95 2.45 14.65 4.60 ;
        RECT  14.25 7.70 14.95 10.55 ;
        RECT  8.85 10.05 14.95 10.55 ;
        RECT  10.20 6.75 16.30 7.25 ;
        RECT  15.60 6.75 16.30 10.55 ;
        RECT  16.65 2.45 17.35 4.60 ;
        RECT  0.45 4.10 17.35 4.60 ;
        RECT  18.00 3.40 18.70 4.10 ;
        RECT  18.30 7.70 19.00 10.55 ;
        RECT  19.35 2.45 20.05 3.15 ;
        RECT  20.70 3.40 21.40 4.10 ;
        RECT  21.00 7.70 21.70 10.55 ;
        RECT  15.60 10.05 21.70 10.55 ;
        RECT  16.65 2.45 22.75 2.95 ;
        RECT  22.05 2.45 22.75 3.15 ;
        RECT  23.60 2.45 24.30 4.10 ;
        RECT  18.00 3.60 24.30 4.10 ;
        RECT  26.30 2.45 27.00 3.15 ;
        RECT  23.60 2.45 29.70 2.95 ;
        RECT  29.00 2.45 29.70 4.10 ;
    END
END ON311X4
MACRO ON31X1
    CLASS CORE ;
    FOREIGN ON31X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.70 6.75 5.20 9.25 ;
        RECT  4.50 7.65 5.20 9.25 ;
        RECT  6.00 2.95 6.50 7.25 ;
        RECT  4.70 6.75 6.50 7.25 ;
        RECT  5.85 2.95 6.55 5.00 ;
        RECT  5.85 4.10 6.75 5.00 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.55 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  3.05 4.10 4.20 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.25 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.75 7.15 1.45 11.00 ;
        RECT  5.85 7.70 6.55 11.00 ;
        RECT  0.00 11.00 7.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.20 3.60 ;
        RECT  3.15 2.00 3.85 2.70 ;
        RECT  0.00 0.00 7.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 2.70 2.50 3.65 ;
        RECT  4.50 2.75 5.20 3.65 ;
        RECT  1.80 3.15 5.20 3.65 ;
    END
END ON31X1
MACRO ON31X2
    CLASS CORE ;
    FOREIGN ON31X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.00 7.70 10.70 10.55 ;
        RECT  12.70 7.15 13.40 10.55 ;
        RECT  12.85 3.40 13.40 10.55 ;
        RECT  10.00 10.05 13.40 10.55 ;
        RECT  12.85 3.40 13.55 4.10 ;
        RECT  12.85 5.40 13.75 6.30 ;
        RECT  12.85 6.75 16.25 7.25 ;
        RECT  12.70 7.15 16.25 7.25 ;
        RECT  15.55 3.40 16.25 4.10 ;
        RECT  12.85 3.60 16.25 4.10 ;
        RECT  15.55 6.75 16.25 10.50 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.80 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.30 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.60 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 11.00 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.60 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.60 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.55 6.75 1.25 11.00 ;
        RECT  0.55 6.75 3.95 7.25 ;
        RECT  3.25 6.75 3.95 9.60 ;
        RECT  14.20 7.70 14.90 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.60 4.10 ;
        RECT  2.65 2.00 3.35 4.00 ;
        RECT  5.35 2.00 6.05 4.00 ;
        RECT  8.05 2.00 8.75 4.00 ;
        RECT  10.75 2.00 11.45 4.00 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.90 7.70 2.60 10.55 ;
        RECT  4.00 2.45 4.70 4.95 ;
        RECT  4.60 6.75 5.30 10.55 ;
        RECT  1.90 10.05 5.30 10.55 ;
        RECT  5.95 7.70 6.65 10.55 ;
        RECT  4.60 6.75 8.00 7.25 ;
        RECT  6.70 2.45 7.40 4.95 ;
        RECT  7.30 6.75 8.00 9.60 ;
        RECT  8.65 6.75 9.35 10.55 ;
        RECT  5.95 10.05 9.35 10.55 ;
        RECT  9.40 2.45 10.10 4.95 ;
        RECT  8.65 6.75 12.05 7.25 ;
        RECT  11.35 6.75 12.05 9.60 ;
        RECT  11.90 2.45 12.40 4.95 ;
        RECT  4.00 4.45 12.40 4.95 ;
        RECT  11.90 2.45 14.90 2.95 ;
        RECT  14.20 2.45 14.90 3.15 ;
    END
END ON31X2
MACRO ON31X4
    CLASS CORE ;
    FOREIGN ON31X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 25.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  15.95 6.75 16.65 9.60 ;
        RECT  18.65 6.75 19.35 9.60 ;
        RECT  20.00 3.40 20.70 4.10 ;
        RECT  21.35 3.60 21.75 10.55 ;
        RECT  21.25 3.60 21.75 7.25 ;
        RECT  21.35 5.40 22.05 10.55 ;
        RECT  21.25 5.40 22.15 7.25 ;
        RECT  22.70 3.40 23.40 4.10 ;
        RECT  20.00 3.60 23.40 4.10 ;
        RECT  15.95 6.75 24.75 7.25 ;
        RECT  24.05 6.75 24.75 10.55 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.60 ;
        PORT
        LAYER M1M ;
        RECT  22.65 5.40 23.55 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 11.20 ;
        PORT
        LAYER M1M ;
        RECT  17.00 5.40 17.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 11.20 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.35 10.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 11.20 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.10 7.15 1.80 11.00 ;
        RECT  3.80 7.70 4.50 11.00 ;
        RECT  6.50 7.70 7.20 11.00 ;
        RECT  22.70 7.70 23.40 11.00 ;
        RECT  0.00 11.00 25.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.70 2.00 1.40 3.80 ;
        RECT  3.80 2.00 4.50 3.65 ;
        RECT  6.50 2.00 7.20 3.65 ;
        RECT  9.20 2.00 9.90 3.65 ;
        RECT  11.90 2.00 12.60 3.65 ;
        RECT  14.60 2.00 15.30 3.65 ;
        RECT  17.30 2.00 18.00 3.65 ;
        RECT  0.00 0.00 25.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.45 2.45 3.15 4.60 ;
        RECT  2.45 6.75 3.15 10.55 ;
        RECT  5.15 2.45 5.85 4.60 ;
        RECT  5.15 6.75 5.85 10.55 ;
        RECT  2.45 6.75 8.55 7.25 ;
        RECT  7.85 2.45 8.55 4.60 ;
        RECT  7.85 6.75 8.55 10.55 ;
        RECT  9.20 6.75 9.90 9.60 ;
        RECT  10.55 2.45 11.25 4.60 ;
        RECT  10.55 7.70 11.25 10.55 ;
        RECT  11.90 6.75 12.60 9.60 ;
        RECT  13.25 2.45 13.95 4.60 ;
        RECT  13.25 7.70 13.95 10.55 ;
        RECT  7.85 10.05 13.95 10.55 ;
        RECT  9.20 6.75 15.30 7.25 ;
        RECT  14.60 6.75 15.30 10.55 ;
        RECT  15.95 2.45 16.65 4.60 ;
        RECT  17.30 7.70 18.00 10.55 ;
        RECT  18.65 2.45 19.35 4.60 ;
        RECT  2.45 4.10 19.35 4.60 ;
        RECT  20.00 7.70 20.70 10.55 ;
        RECT  14.60 10.05 20.70 10.55 ;
        RECT  21.35 2.45 22.05 3.15 ;
        RECT  18.65 2.45 24.75 2.95 ;
        RECT  24.05 2.45 24.75 3.15 ;
    END
END ON31X4
MACRO ON321X1
    CLASS CORE ;
    FOREIGN ON321X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.45 1.15 4.50 ;
        RECT  0.25 5.40 1.15 6.30 ;
        RECT  0.65 2.45 1.15 7.25 ;
        RECT  1.70 6.75 2.40 9.10 ;
        RECT  0.65 6.75 6.10 7.25 ;
        RECT  5.60 6.75 6.10 10.55 ;
        RECT  5.60 7.40 6.30 10.55 ;
        RECT  5.60 7.40 7.40 8.10 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.60 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  5.15 5.40 6.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  7.20 5.40 8.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  8.60 5.25 9.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 10.10 2.35 11.00 ;
        RECT  3.20 7.70 3.90 11.00 ;
        RECT  10.05 7.15 10.75 11.00 ;
        RECT  8.95 10.75 10.75 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  7.35 2.00 8.05 3.45 ;
        RECT  10.05 2.00 10.75 4.10 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 2.45 2.50 4.50 ;
        RECT  3.30 3.70 4.00 4.40 ;
        RECT  1.80 2.45 5.35 2.95 ;
        RECT  4.65 2.45 5.35 3.40 ;
        RECT  6.00 2.45 6.70 4.40 ;
        RECT  8.70 2.45 9.40 4.40 ;
        RECT  3.30 3.90 9.40 4.40 ;
    END
END ON321X1
MACRO ON321X2
    CLASS CORE ;
    FOREIGN ON321X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  2.60 7.10 3.30 10.55 ;
        RECT  0.45 3.80 3.95 4.50 ;
        RECT  3.05 5.40 3.95 6.30 ;
        RECT  3.45 3.80 3.95 7.60 ;
        RECT  2.60 7.10 6.80 7.60 ;
        RECT  6.30 7.10 6.80 8.55 ;
        RECT  6.30 7.85 10.10 8.55 ;
        RECT  6.30 8.05 17.20 8.55 ;
        RECT  9.40 7.85 10.10 10.55 ;
        RECT  16.50 7.15 17.20 8.75 ;
        RECT  9.40 8.05 17.20 8.75 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.50 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.60 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  10.00 5.40 10.95 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  4.40 5.40 5.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  14.20 5.40 15.15 6.35 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  18.15 5.25 19.35 5.95 ;
        RECT  18.45 5.25 19.35 6.35 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.75 9.55 1.45 11.00 ;
        RECT  3.95 8.05 4.65 11.00 ;
        RECT  3.95 10.20 7.75 11.00 ;
        RECT  19.85 7.15 20.55 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  11.95 2.00 12.65 3.55 ;
        RECT  14.65 2.00 15.35 3.55 ;
        RECT  14.65 2.85 17.85 3.55 ;
        RECT  19.85 2.00 20.55 4.50 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.45 2.45 4.30 3.15 ;
        RECT  5.95 3.80 8.80 4.50 ;
        RECT  6.95 2.45 9.80 3.15 ;
        RECT  1.45 2.65 9.80 3.15 ;
        RECT  10.45 2.45 11.15 4.50 ;
        RECT  13.30 2.45 14.00 4.50 ;
        RECT  18.50 2.55 19.20 4.50 ;
        RECT  5.95 4.00 19.20 4.50 ;
    END
END ON321X2
MACRO ON321X4
    CLASS CORE ;
    FOREIGN ON321X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 39.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  16.95 6.75 17.65 9.60 ;
        RECT  19.65 6.75 20.35 9.60 ;
        RECT  22.35 6.75 23.05 10.55 ;
        RECT  25.05 8.65 25.75 10.55 ;
        RECT  27.75 8.65 28.45 10.55 ;
        RECT  22.35 10.05 28.45 10.55 ;
        RECT  32.45 3.40 32.95 7.25 ;
        RECT  32.45 3.40 33.20 4.10 ;
        RECT  32.45 5.40 33.35 7.25 ;
        RECT  35.20 3.40 35.90 4.10 ;
        RECT  32.45 3.60 35.90 4.10 ;
        RECT  16.95 6.75 36.70 7.25 ;
        RECT  36.00 6.75 36.70 10.55 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 7.00 ;
        PORT
        LAYER M1M ;
        RECT  35.25 5.40 36.15 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  22.65 5.40 23.55 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  29.65 5.40 30.55 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.55 9.60 1.25 11.00 ;
        RECT  2.10 7.15 2.80 11.00 ;
        RECT  4.80 7.70 5.50 11.00 ;
        RECT  7.50 7.70 8.20 11.00 ;
        RECT  29.25 8.65 29.95 11.00 ;
        RECT  31.95 8.65 32.65 11.00 ;
        RECT  34.65 7.70 35.35 11.00 ;
        RECT  37.35 7.10 38.05 11.00 ;
        RECT  0.00 11.00 39.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.55 2.00 1.25 4.25 ;
        RECT  4.00 2.00 4.70 3.60 ;
        RECT  6.70 2.00 7.40 3.60 ;
        RECT  9.40 2.00 10.10 3.60 ;
        RECT  12.10 2.00 12.80 3.60 ;
        RECT  14.80 2.00 15.50 3.60 ;
        RECT  17.50 2.00 18.20 3.60 ;
        RECT  38.05 2.00 38.75 4.10 ;
        RECT  0.00 0.00 39.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.65 2.45 3.35 4.60 ;
        RECT  3.45 6.75 4.15 10.55 ;
        RECT  5.35 2.45 6.05 4.60 ;
        RECT  6.15 6.75 6.85 10.55 ;
        RECT  8.05 2.45 8.75 4.60 ;
        RECT  3.45 6.75 9.55 7.25 ;
        RECT  8.85 6.75 9.55 10.55 ;
        RECT  10.20 6.75 10.90 9.60 ;
        RECT  10.75 2.45 11.45 4.60 ;
        RECT  11.55 7.70 12.25 10.55 ;
        RECT  12.90 6.75 13.60 9.60 ;
        RECT  13.45 2.45 14.15 4.60 ;
        RECT  14.25 7.70 14.95 10.55 ;
        RECT  8.85 10.05 14.95 10.55 ;
        RECT  10.20 6.75 16.30 7.25 ;
        RECT  15.60 6.75 16.30 10.55 ;
        RECT  16.15 2.45 16.85 4.60 ;
        RECT  18.30 7.70 19.00 10.55 ;
        RECT  18.85 2.45 19.55 4.60 ;
        RECT  2.65 4.10 19.55 4.60 ;
        RECT  20.20 3.40 20.90 4.10 ;
        RECT  21.00 7.70 21.70 10.55 ;
        RECT  15.60 10.05 21.70 10.55 ;
        RECT  21.55 2.45 22.25 3.15 ;
        RECT  22.90 3.40 23.60 4.10 ;
        RECT  23.70 7.70 24.40 9.60 ;
        RECT  24.25 2.45 24.95 3.15 ;
        RECT  25.60 3.40 26.30 4.10 ;
        RECT  26.40 7.70 27.10 9.60 ;
        RECT  26.95 2.45 27.65 3.15 ;
        RECT  28.30 3.40 29.00 4.10 ;
        RECT  18.85 2.45 30.35 2.95 ;
        RECT  29.65 2.45 30.35 3.15 ;
        RECT  30.60 7.70 31.30 10.55 ;
        RECT  31.15 2.45 31.85 4.10 ;
        RECT  20.20 3.60 31.85 4.10 ;
        RECT  23.70 7.70 34.00 8.20 ;
        RECT  33.30 7.70 34.00 10.55 ;
        RECT  33.85 2.45 34.55 3.15 ;
        RECT  31.15 2.45 37.25 2.95 ;
        RECT  36.55 2.45 37.25 4.10 ;
    END
END ON321X4
MACRO ON322X1
    CLASS CORE ;
    FOREIGN ON322X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  3.80 7.20 4.50 8.80 ;
        RECT  4.90 8.30 5.60 10.55 ;
        RECT  7.45 6.85 7.95 8.80 ;
        RECT  3.80 8.30 7.95 8.80 ;
        RECT  10.05 3.55 10.55 7.35 ;
        RECT  10.05 3.55 10.80 4.25 ;
        RECT  10.05 5.40 10.95 6.30 ;
        RECT  7.45 6.85 12.15 7.35 ;
        RECT  11.45 6.85 12.15 10.55 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.40 9.55 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  5.85 6.70 6.75 7.60 ;
        RECT  5.40 6.85 6.75 7.60 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  4.15 5.40 5.35 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.35 2.90 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.15 1.15 11.00 ;
        RECT  7.25 9.25 7.95 11.00 ;
        RECT  9.10 7.85 9.80 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 4.45 ;
        RECT  3.10 2.00 3.90 3.30 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 2.55 2.50 4.25 ;
        RECT  4.50 2.45 5.20 4.25 ;
        RECT  1.80 3.75 5.20 4.25 ;
        RECT  5.85 3.70 6.55 4.40 ;
        RECT  4.50 2.45 7.90 2.95 ;
        RECT  7.20 2.45 7.90 3.15 ;
        RECT  8.75 2.55 9.45 4.40 ;
        RECT  5.85 3.90 9.45 4.40 ;
        RECT  8.75 2.55 12.15 3.05 ;
        RECT  11.45 2.55 12.15 4.40 ;
    END
END ON322X1
MACRO ON322X2
    CLASS CORE ;
    FOREIGN ON322X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  3.80 7.15 4.50 8.75 ;
        RECT  3.80 8.05 11.60 8.75 ;
        RECT  10.90 7.85 11.60 10.55 ;
        RECT  10.90 7.85 14.70 8.55 ;
        RECT  14.20 7.10 14.70 8.55 ;
        RECT  3.80 8.05 14.70 8.55 ;
        RECT  14.20 7.10 19.20 7.60 ;
        RECT  18.70 7.10 19.20 8.55 ;
        RECT  16.85 3.80 22.20 4.50 ;
        RECT  21.25 5.40 22.20 6.30 ;
        RECT  18.70 7.85 22.50 8.55 ;
        RECT  21.80 3.80 22.20 10.55 ;
        RECT  21.70 3.80 22.20 8.55 ;
        RECT  21.80 7.85 22.50 10.55 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.30 17.95 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.35 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.80 6.35 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.35 2.90 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.15 1.15 11.00 ;
        RECT  16.35 8.05 17.05 11.00 ;
        RECT  13.25 10.20 20.15 11.00 ;
        RECT  0.00 11.00 23.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 4.50 ;
        RECT  5.65 2.00 6.35 3.55 ;
        RECT  3.15 2.85 6.35 3.55 ;
        RECT  8.35 2.00 9.05 3.55 ;
        RECT  0.00 0.00 23.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 2.55 2.50 4.50 ;
        RECT  7.00 2.45 7.70 4.50 ;
        RECT  9.85 2.45 10.55 4.50 ;
        RECT  11.20 2.45 14.05 3.15 ;
        RECT  12.20 3.80 15.05 4.50 ;
        RECT  1.80 4.00 15.05 4.50 ;
        RECT  15.85 2.45 18.70 3.15 ;
        RECT  20.35 2.45 23.20 3.15 ;
        RECT  11.20 2.65 23.20 3.15 ;
    END
END ON322X2
MACRO ON322X4
    CLASS CORE ;
    FOREIGN ON322X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 49.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  16.95 6.75 17.65 9.60 ;
        RECT  19.65 6.75 20.35 9.60 ;
        RECT  22.35 6.75 23.05 10.55 ;
        RECT  25.05 8.65 25.75 10.55 ;
        RECT  27.75 8.65 28.45 10.55 ;
        RECT  22.35 10.05 28.45 10.55 ;
        RECT  34.50 3.40 35.20 4.10 ;
        RECT  37.20 3.40 37.90 4.10 ;
        RECT  38.05 3.60 38.55 7.25 ;
        RECT  38.05 5.40 38.95 7.25 ;
        RECT  39.90 3.40 40.60 4.10 ;
        RECT  42.60 3.40 43.30 4.10 ;
        RECT  34.50 3.60 43.30 4.10 ;
        RECT  42.90 6.75 43.60 9.60 ;
        RECT  16.95 6.75 46.30 7.25 ;
        RECT  45.60 6.75 46.30 9.60 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  42.25 5.40 43.15 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  35.25 5.40 36.15 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  22.65 5.40 23.55 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  29.65 5.40 30.55 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.55 9.60 1.25 11.00 ;
        RECT  2.10 7.15 2.80 11.00 ;
        RECT  4.80 7.70 5.50 11.00 ;
        RECT  7.50 7.70 8.20 11.00 ;
        RECT  29.25 8.65 29.95 11.00 ;
        RECT  31.95 8.65 32.65 11.00 ;
        RECT  34.65 7.70 35.35 11.00 ;
        RECT  37.35 8.65 38.05 11.00 ;
        RECT  40.05 8.65 40.75 11.00 ;
        RECT  0.00 11.00 49.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 3.85 4.25 ;
        RECT  6.00 2.00 6.70 3.60 ;
        RECT  8.70 2.00 9.40 3.60 ;
        RECT  11.40 2.00 12.10 3.60 ;
        RECT  14.10 2.00 14.80 3.60 ;
        RECT  16.80 2.00 17.50 3.60 ;
        RECT  19.50 2.00 20.20 3.60 ;
        RECT  45.45 2.00 48.55 4.25 ;
        RECT  0.00 0.00 49.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.45 6.75 4.15 10.55 ;
        RECT  4.65 2.45 5.35 4.60 ;
        RECT  6.15 6.75 6.85 10.55 ;
        RECT  7.35 2.45 8.05 4.60 ;
        RECT  3.45 6.75 9.55 7.25 ;
        RECT  8.85 6.75 9.55 10.55 ;
        RECT  10.05 2.45 10.75 4.60 ;
        RECT  10.20 6.75 10.90 9.60 ;
        RECT  11.55 7.70 12.25 10.55 ;
        RECT  12.75 2.45 13.45 4.60 ;
        RECT  12.90 6.75 13.60 9.60 ;
        RECT  14.25 7.70 14.95 10.55 ;
        RECT  8.85 10.05 14.95 10.55 ;
        RECT  10.20 6.75 16.30 7.25 ;
        RECT  15.45 2.45 16.15 4.60 ;
        RECT  15.60 6.75 16.30 10.55 ;
        RECT  18.15 2.45 18.85 4.60 ;
        RECT  18.30 7.70 19.00 10.55 ;
        RECT  20.85 2.45 21.55 4.60 ;
        RECT  4.65 4.10 21.55 4.60 ;
        RECT  21.00 7.70 21.70 10.55 ;
        RECT  15.60 10.05 21.70 10.55 ;
        RECT  22.20 3.40 22.90 4.10 ;
        RECT  23.55 2.45 24.25 3.15 ;
        RECT  23.70 7.70 24.40 9.60 ;
        RECT  24.90 3.40 25.60 4.10 ;
        RECT  26.25 2.45 26.95 3.15 ;
        RECT  26.40 7.70 27.10 9.60 ;
        RECT  27.60 3.40 28.30 4.10 ;
        RECT  28.95 2.45 29.65 3.15 ;
        RECT  30.30 3.40 31.00 4.10 ;
        RECT  30.60 7.70 31.30 10.55 ;
        RECT  20.85 2.45 32.35 2.95 ;
        RECT  31.65 2.45 32.35 3.15 ;
        RECT  23.70 7.70 34.00 8.20 ;
        RECT  33.15 2.45 33.85 4.10 ;
        RECT  22.20 3.60 33.85 4.10 ;
        RECT  33.30 7.70 34.00 10.55 ;
        RECT  35.85 2.45 36.55 3.15 ;
        RECT  36.00 7.70 36.70 10.55 ;
        RECT  38.55 2.45 39.25 3.15 ;
        RECT  38.70 7.70 39.40 10.55 ;
        RECT  36.00 7.70 42.25 8.20 ;
        RECT  41.25 2.45 41.95 3.15 ;
        RECT  41.55 7.70 42.25 10.55 ;
        RECT  33.15 2.45 44.65 2.95 ;
        RECT  43.95 2.45 44.65 4.10 ;
        RECT  44.25 7.70 44.95 10.55 ;
        RECT  46.95 7.70 47.65 10.55 ;
        RECT  41.55 10.05 47.65 10.55 ;
    END
END ON322X4
MACRO ON32X1
    CLASS CORE ;
    FOREIGN ON32X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  3.80 7.10 5.55 7.80 ;
        RECT  4.85 7.10 5.55 10.55 ;
        RECT  5.85 3.40 6.35 7.65 ;
        RECT  3.80 7.10 6.35 7.65 ;
        RECT  5.85 3.40 6.55 4.10 ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.25 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.15 1.15 11.00 ;
        RECT  0.45 10.45 2.20 11.00 ;
        RECT  7.20 7.25 7.90 11.00 ;
        RECT  0.00 11.00 8.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.20 3.90 ;
        RECT  3.15 2.00 3.85 3.00 ;
        RECT  0.00 0.00 8.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 2.45 2.50 4.05 ;
        RECT  4.50 2.45 5.20 4.05 ;
        RECT  1.80 3.55 5.20 4.05 ;
        RECT  4.50 2.45 7.90 2.95 ;
        RECT  7.20 2.45 7.90 4.05 ;
    END
END ON32X1
MACRO ON32X2
    CLASS CORE ;
    FOREIGN ON32X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.00 7.70 10.70 10.55 ;
        RECT  12.85 3.40 13.40 10.55 ;
        RECT  12.70 7.15 13.40 10.55 ;
        RECT  12.85 3.40 13.55 4.95 ;
        RECT  12.85 5.40 13.75 6.30 ;
        RECT  15.40 7.70 16.10 10.55 ;
        RECT  10.00 10.05 16.10 10.55 ;
        RECT  15.55 3.40 16.25 4.95 ;
        RECT  18.25 2.45 18.95 4.95 ;
        RECT  12.85 4.45 18.95 4.95 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.20 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.20 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.20 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 18.00 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.60 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 11.00 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.60 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.60 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.55 6.75 1.25 11.00 ;
        RECT  0.55 6.75 3.95 7.25 ;
        RECT  3.25 6.75 3.95 9.60 ;
        RECT  16.90 7.70 17.60 11.00 ;
        RECT  19.60 7.70 20.30 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.65 2.00 1.35 4.00 ;
        RECT  2.65 2.00 3.35 4.00 ;
        RECT  5.35 2.00 6.05 4.00 ;
        RECT  8.05 2.00 8.75 4.00 ;
        RECT  10.75 2.00 11.45 4.00 ;
        RECT  19.75 2.00 20.45 4.00 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.90 7.70 2.60 10.55 ;
        RECT  4.00 2.45 4.70 4.95 ;
        RECT  4.60 6.75 5.30 10.55 ;
        RECT  1.90 10.05 5.30 10.55 ;
        RECT  5.95 7.70 6.65 10.55 ;
        RECT  4.60 6.75 8.00 7.25 ;
        RECT  6.70 2.45 7.40 4.95 ;
        RECT  7.30 6.75 8.00 9.60 ;
        RECT  8.65 6.75 9.35 10.55 ;
        RECT  5.95 10.05 9.35 10.55 ;
        RECT  9.40 2.45 10.10 4.95 ;
        RECT  8.65 6.75 12.05 7.25 ;
        RECT  11.35 6.75 12.05 9.60 ;
        RECT  11.90 2.45 12.40 4.95 ;
        RECT  4.00 4.45 12.40 4.95 ;
        RECT  14.05 6.75 14.75 9.60 ;
        RECT  14.20 2.45 14.90 3.15 ;
        RECT  11.90 2.45 17.60 2.95 ;
        RECT  16.90 2.45 17.60 3.15 ;
        RECT  14.05 6.75 18.95 7.25 ;
        RECT  18.25 6.75 18.95 10.50 ;
    END
END ON32X2
MACRO ON32X4
    CLASS CORE ;
    FOREIGN ON32X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 30.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  15.30 6.75 16.00 9.60 ;
        RECT  18.00 6.75 18.70 9.60 ;
        RECT  15.30 6.75 21.40 7.25 ;
        RECT  20.20 3.40 20.75 7.25 ;
        RECT  20.70 3.40 20.75 10.55 ;
        RECT  19.85 5.40 20.75 7.25 ;
        RECT  20.20 3.40 20.90 4.10 ;
        RECT  20.70 6.75 21.40 10.55 ;
        RECT  22.90 3.40 23.60 4.10 ;
        RECT  25.60 3.40 26.30 4.10 ;
        RECT  20.70 9.15 27.05 9.85 ;
        RECT  28.30 3.40 29.00 4.10 ;
        RECT  20.20 3.60 29.00 4.10 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 8.40 ;
        PORT
        LAYER M1M ;
        RECT  21.25 5.40 22.15 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 8.40 ;
        PORT
        LAYER M1M ;
        RECT  24.05 5.40 24.95 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 11.20 ;
        PORT
        LAYER M1M ;
        RECT  17.00 5.35 17.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 11.20 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.35 10.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 11.20 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.15 1.15 11.00 ;
        RECT  3.15 7.70 3.85 11.00 ;
        RECT  5.85 7.70 6.55 11.00 ;
        RECT  23.20 6.80 29.40 7.50 ;
        RECT  28.70 6.80 29.40 11.00 ;
        RECT  0.00 11.00 30.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.80 2.00 1.50 3.80 ;
        RECT  4.00 2.00 4.70 3.65 ;
        RECT  6.70 2.00 7.40 3.65 ;
        RECT  9.40 2.00 10.10 3.65 ;
        RECT  12.10 2.00 12.80 3.65 ;
        RECT  14.80 2.00 15.50 3.65 ;
        RECT  17.50 2.00 18.20 3.65 ;
        RECT  0.00 0.00 30.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 6.75 2.50 10.55 ;
        RECT  2.65 2.45 3.35 4.60 ;
        RECT  4.50 6.75 5.20 10.55 ;
        RECT  5.35 2.45 6.05 4.60 ;
        RECT  1.80 6.75 7.90 7.25 ;
        RECT  7.20 6.75 7.90 10.55 ;
        RECT  8.05 2.45 8.75 4.60 ;
        RECT  8.55 6.75 9.25 9.60 ;
        RECT  9.90 7.70 10.60 10.55 ;
        RECT  10.75 2.45 11.45 4.60 ;
        RECT  11.25 6.75 11.95 9.60 ;
        RECT  12.60 7.70 13.30 10.55 ;
        RECT  7.20 10.05 13.30 10.55 ;
        RECT  8.55 6.75 14.65 7.25 ;
        RECT  13.45 2.45 14.15 4.60 ;
        RECT  13.95 6.75 14.65 10.55 ;
        RECT  16.15 2.45 16.85 4.60 ;
        RECT  16.65 7.70 17.35 10.55 ;
        RECT  18.85 2.45 19.55 4.60 ;
        RECT  2.65 4.10 19.55 4.60 ;
        RECT  19.35 7.70 20.05 10.55 ;
        RECT  13.95 10.05 20.05 10.55 ;
        RECT  21.55 2.45 22.25 3.15 ;
        RECT  24.25 2.45 24.95 3.15 ;
        RECT  26.95 2.45 27.65 3.15 ;
        RECT  18.85 2.45 30.35 2.95 ;
        RECT  29.65 2.45 30.35 3.15 ;
    END
END ON32X4
MACRO ON331X1
    CLASS CORE ;
    FOREIGN ON331X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        RECT  1.05 4.30 1.15 8.80 ;
        RECT  0.65 4.30 1.15 7.65 ;
        RECT  1.05 7.15 1.75 8.80 ;
        RECT  1.95 2.55 2.65 4.80 ;
        RECT  0.65 4.30 2.65 4.80 ;
        RECT  0.65 7.15 6.40 7.65 ;
        RECT  5.90 7.15 6.40 8.85 ;
        RECT  7.00 8.05 7.70 10.55 ;
        RECT  5.90 8.05 8.80 8.85 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.35 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.35 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.35 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.35 8.90 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  9.60 5.40 10.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.15 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.70 10.10 1.40 11.00 ;
        RECT  2.55 8.35 3.25 11.00 ;
        RECT  11.45 7.15 12.15 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.80 ;
        RECT  8.70 2.00 9.40 3.30 ;
        RECT  11.40 2.00 12.10 4.45 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.30 2.55 4.00 4.35 ;
        RECT  4.65 3.55 5.35 4.25 ;
        RECT  3.30 2.55 6.70 3.05 ;
        RECT  6.00 2.55 6.70 3.25 ;
        RECT  7.35 2.55 8.05 4.25 ;
        RECT  10.05 2.55 10.75 4.25 ;
        RECT  4.65 3.75 10.75 4.25 ;
    END
END ON331X1
MACRO ON331X2
    CLASS CORE ;
    FOREIGN ON331X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 25.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.45 0.75 10.55 ;
        RECT  0.25 2.45 0.75 7.65 ;
        RECT  0.25 5.40 1.15 6.30 ;
        RECT  0.45 7.15 1.20 10.55 ;
        RECT  0.25 2.45 3.35 3.15 ;
        RECT  0.25 7.15 6.05 7.65 ;
        RECT  5.55 7.15 6.05 8.80 ;
        RECT  12.45 8.05 13.15 10.55 ;
        RECT  19.55 7.15 20.25 8.80 ;
        RECT  5.55 8.05 20.25 8.80 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.50 ;
        PORT
        LAYER M1M ;
        RECT  1.60 5.40 2.55 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.25 10.95 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.25 3.95 6.35 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.40 19.45 6.35 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.28 ;
        PORT
        LAYER M1M ;
        RECT  21.25 5.35 22.15 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.28 ;
        PORT
        LAYER M1M ;
        RECT  22.60 5.40 23.55 6.35 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.00 8.10 2.70 11.00 ;
        RECT  22.90 7.10 23.60 11.00 ;
        RECT  0.00 11.00 25.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  16.20 2.00 16.90 3.55 ;
        RECT  18.90 2.00 19.60 3.55 ;
        RECT  18.90 2.85 22.05 3.55 ;
        RECT  24.05 2.00 24.75 4.45 ;
        RECT  0.00 0.00 25.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.95 2.45 4.45 4.50 ;
        RECT  1.50 3.80 4.45 4.50 ;
        RECT  3.95 2.45 13.90 3.15 ;
        RECT  14.55 2.45 15.25 4.50 ;
        RECT  5.05 3.80 15.25 4.50 ;
        RECT  17.55 2.45 18.25 4.50 ;
        RECT  22.70 2.55 23.40 4.50 ;
        RECT  5.05 4.00 23.40 4.50 ;
    END
END ON331X2
MACRO ON331X4
    CLASS CORE ;
    FOREIGN ON331X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 50.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  16.95 6.75 17.65 9.60 ;
        RECT  19.65 6.75 20.35 9.60 ;
        RECT  22.35 6.75 23.05 10.55 ;
        RECT  32.40 5.80 32.90 7.25 ;
        RECT  16.95 6.75 32.90 7.25 ;
        RECT  32.40 5.80 40.40 6.30 ;
        RECT  40.20 5.80 40.40 9.60 ;
        RECT  39.90 5.80 40.40 7.25 ;
        RECT  40.20 6.75 40.90 9.60 ;
        RECT  42.90 6.75 43.60 9.60 ;
        RECT  43.80 3.40 44.55 4.10 ;
        RECT  44.05 3.40 44.55 7.25 ;
        RECT  43.65 5.40 44.55 7.25 ;
        RECT  45.60 6.75 46.30 10.55 ;
        RECT  46.50 3.40 47.20 4.10 ;
        RECT  39.90 6.75 49.00 7.25 ;
        RECT  48.30 6.75 49.00 10.55 ;
        RECT  49.20 2.45 49.90 4.10 ;
        RECT  43.80 3.60 49.90 4.10 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 7.00 ;
        PORT
        LAYER M1M ;
        RECT  46.45 5.40 47.35 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  40.85 5.40 41.75 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  31.05 5.40 31.95 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  26.85 5.40 27.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.40 19.35 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.55 9.55 1.25 11.00 ;
        RECT  2.10 7.15 2.80 11.00 ;
        RECT  4.80 7.70 5.50 11.00 ;
        RECT  7.50 7.70 8.20 11.00 ;
        RECT  23.85 7.70 24.55 11.00 ;
        RECT  25.35 7.70 26.05 11.00 ;
        RECT  28.05 8.65 28.75 11.00 ;
        RECT  30.75 8.70 31.45 11.00 ;
        RECT  46.95 7.70 47.65 11.00 ;
        RECT  0.00 11.00 50.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 4.25 ;
        RECT  1.95 2.00 2.65 3.80 ;
        RECT  4.65 2.00 5.35 3.80 ;
        RECT  7.35 2.00 8.05 3.80 ;
        RECT  10.05 2.00 10.75 3.80 ;
        RECT  12.75 2.00 13.45 3.80 ;
        RECT  15.45 2.00 16.15 3.80 ;
        RECT  18.15 2.00 18.85 3.80 ;
        RECT  20.85 2.00 21.55 3.80 ;
        RECT  0.00 0.00 50.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.30 2.45 4.00 4.80 ;
        RECT  3.45 6.75 4.15 10.55 ;
        RECT  6.00 2.45 6.70 4.80 ;
        RECT  6.15 6.75 6.85 10.55 ;
        RECT  3.45 6.75 9.55 7.25 ;
        RECT  8.70 2.45 9.40 4.80 ;
        RECT  8.85 6.75 9.55 10.55 ;
        RECT  10.20 6.75 10.90 9.60 ;
        RECT  11.40 2.45 12.10 4.80 ;
        RECT  11.55 7.70 12.25 10.55 ;
        RECT  12.90 6.75 13.60 9.60 ;
        RECT  14.10 2.45 14.80 4.80 ;
        RECT  14.25 7.70 14.95 10.55 ;
        RECT  8.85 10.05 14.95 10.55 ;
        RECT  10.20 6.75 16.30 7.25 ;
        RECT  15.60 6.75 16.30 10.55 ;
        RECT  16.80 2.45 17.50 4.80 ;
        RECT  18.30 7.70 19.00 10.55 ;
        RECT  19.50 2.45 20.20 4.80 ;
        RECT  21.00 7.70 21.70 10.55 ;
        RECT  15.60 10.05 21.70 10.55 ;
        RECT  22.20 2.45 22.90 4.80 ;
        RECT  3.30 4.30 22.90 4.80 ;
        RECT  23.55 3.40 24.25 4.10 ;
        RECT  24.90 2.45 25.60 3.15 ;
        RECT  26.25 3.40 26.95 4.10 ;
        RECT  26.70 7.70 27.40 10.55 ;
        RECT  27.60 2.45 28.30 3.15 ;
        RECT  28.95 3.40 29.65 4.10 ;
        RECT  29.40 7.70 30.10 10.55 ;
        RECT  30.30 2.45 31.00 3.15 ;
        RECT  26.70 7.70 32.80 8.20 ;
        RECT  31.65 3.40 32.35 4.10 ;
        RECT  32.10 7.70 32.80 10.55 ;
        RECT  33.00 2.45 33.70 3.15 ;
        RECT  33.45 6.75 34.15 9.60 ;
        RECT  34.35 3.40 35.05 4.10 ;
        RECT  34.80 7.70 35.50 10.55 ;
        RECT  35.70 2.45 36.40 3.15 ;
        RECT  36.15 6.75 36.85 9.60 ;
        RECT  37.05 3.40 37.75 4.10 ;
        RECT  37.50 7.70 38.20 10.55 ;
        RECT  32.10 10.05 38.20 10.55 ;
        RECT  33.45 6.75 39.35 7.25 ;
        RECT  38.40 2.45 39.10 3.15 ;
        RECT  38.85 6.75 39.35 10.55 ;
        RECT  38.85 7.70 39.55 10.55 ;
        RECT  39.75 3.40 40.45 4.10 ;
        RECT  22.20 2.45 41.80 2.95 ;
        RECT  41.10 2.45 41.80 3.15 ;
        RECT  41.55 7.70 42.25 10.55 ;
        RECT  42.45 2.45 43.15 4.10 ;
        RECT  23.55 3.60 43.15 4.10 ;
        RECT  44.25 7.70 44.95 10.55 ;
        RECT  38.85 10.05 44.95 10.55 ;
        RECT  45.15 2.45 45.85 3.15 ;
        RECT  42.45 2.45 48.55 2.95 ;
        RECT  47.85 2.45 48.55 3.15 ;
    END
END ON331X4
MACRO ON332X1
    CLASS CORE ;
    FOREIGN ON332X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        RECT  0.65 3.75 1.15 10.00 ;
        RECT  0.45 7.20 1.15 10.00 ;
        RECT  2.05 6.90 2.55 7.90 ;
        RECT  0.45 7.20 2.55 7.90 ;
        RECT  3.40 3.55 4.10 4.25 ;
        RECT  0.65 3.75 4.10 4.25 ;
        RECT  2.05 6.90 6.45 7.40 ;
        RECT  0.45 7.20 6.45 7.40 ;
        RECT  5.95 6.90 6.45 8.55 ;
        RECT  5.95 8.05 10.20 8.55 ;
        RECT  7.40 8.05 9.15 8.85 ;
        RECT  8.45 8.05 9.15 10.55 ;
        RECT  7.40 8.05 10.20 8.80 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 4.00 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.35 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.35 6.75 6.35 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.35 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  9.95 5.40 10.95 6.35 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.25 12.35 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.35 13.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  4.05 7.85 4.75 11.00 ;
        RECT  12.85 7.15 13.55 11.00 ;
        RECT  0.00 11.00 14.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.30 ;
        RECT  10.15 2.00 10.85 3.45 ;
        RECT  12.85 2.00 13.55 3.35 ;
        RECT  0.00 0.00 14.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  2.00 2.55 2.70 3.25 ;
        RECT  4.75 2.55 5.45 3.25 ;
        RECT  6.10 3.55 6.80 4.45 ;
        RECT  2.00 2.55 8.15 3.05 ;
        RECT  7.45 2.55 8.15 3.45 ;
        RECT  8.80 2.55 9.50 4.45 ;
        RECT  11.50 2.55 12.20 4.45 ;
        RECT  6.10 3.95 12.20 4.45 ;
    END
END ON332X1
MACRO ON332X2
    CLASS CORE ;
    FOREIGN ON332X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 30.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  2.15 8.95 2.85 10.55 ;
        RECT  5.25 7.15 5.95 9.70 ;
        RECT  5.85 3.80 5.95 9.70 ;
        RECT  2.15 8.95 5.95 9.70 ;
        RECT  5.85 3.80 6.35 7.65 ;
        RECT  5.85 5.40 6.75 6.30 ;
        RECT  1.80 3.80 7.15 4.50 ;
        RECT  5.25 7.15 11.65 7.65 ;
        RECT  11.15 7.15 11.65 8.80 ;
        RECT  18.05 8.05 18.75 10.55 ;
        RECT  25.15 7.15 25.85 8.80 ;
        RECT  11.15 8.05 25.85 8.80 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  1.55 5.40 2.55 6.30 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.90 ;
        PORT
        LAYER M1M ;
        RECT  7.20 5.40 8.15 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 17.95 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.25 16.55 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.25 9.55 6.35 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  24.05 5.40 25.05 6.35 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.28 ;
        PORT
        LAYER M1M ;
        RECT  26.85 5.35 27.75 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.28 ;
        PORT
        LAYER M1M ;
        RECT  28.20 5.40 29.15 6.35 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.55 9.55 1.25 11.00 ;
        RECT  7.60 8.10 8.30 11.00 ;
        RECT  28.50 7.10 29.20 11.00 ;
        RECT  0.00 11.00 30.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  21.80 2.00 22.50 3.55 ;
        RECT  24.50 2.00 25.20 3.55 ;
        RECT  24.50 2.85 27.65 3.55 ;
        RECT  29.65 2.00 30.35 4.45 ;
        RECT  0.00 0.00 30.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 2.45 1.15 4.50 ;
        RECT  7.80 2.45 8.50 4.50 ;
        RECT  9.30 2.45 10.00 4.50 ;
        RECT  0.45 2.45 19.50 3.15 ;
        RECT  20.15 2.45 20.85 4.50 ;
        RECT  10.65 3.80 20.85 4.50 ;
        RECT  23.15 2.45 23.85 4.50 ;
        RECT  28.30 2.55 29.00 4.50 ;
        RECT  10.65 4.00 29.00 4.50 ;
    END
END ON332X2
MACRO ON332X4
    CLASS CORE ;
    FOREIGN ON332X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 60.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  16.95 6.75 17.65 9.60 ;
        RECT  19.65 6.75 20.35 9.60 ;
        RECT  22.35 6.75 23.05 10.55 ;
        RECT  32.40 5.80 32.90 7.25 ;
        RECT  16.95 6.75 32.90 7.25 ;
        RECT  32.40 5.80 40.40 6.30 ;
        RECT  40.20 5.80 40.40 9.60 ;
        RECT  39.90 5.80 40.40 7.25 ;
        RECT  40.20 6.75 40.90 9.60 ;
        RECT  42.90 6.75 43.60 9.60 ;
        RECT  43.80 3.40 44.55 4.10 ;
        RECT  44.05 3.40 44.55 7.25 ;
        RECT  43.65 5.40 44.55 7.25 ;
        RECT  45.60 6.75 46.30 10.55 ;
        RECT  46.50 3.40 47.20 4.10 ;
        RECT  48.45 6.75 49.15 9.60 ;
        RECT  49.20 3.40 49.90 4.10 ;
        RECT  39.90 6.75 51.85 7.25 ;
        RECT  51.15 6.75 51.85 9.60 ;
        RECT  51.90 3.40 52.60 4.10 ;
        RECT  54.60 3.40 55.30 4.10 ;
        RECT  43.80 3.60 55.30 4.10 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  47.85 5.40 48.75 6.30 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 9.80 ;
        PORT
        LAYER M1M ;
        RECT  53.45 5.40 54.35 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  40.85 5.40 41.75 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  31.05 5.40 31.95 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  26.85 5.40 27.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.40 19.35 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.55 9.55 1.25 11.00 ;
        RECT  2.10 7.15 2.80 11.00 ;
        RECT  4.80 7.70 5.50 11.00 ;
        RECT  7.50 7.70 8.20 11.00 ;
        RECT  23.85 7.70 24.55 11.00 ;
        RECT  25.35 7.70 26.05 11.00 ;
        RECT  28.05 8.65 28.75 11.00 ;
        RECT  30.75 8.70 31.45 11.00 ;
        RECT  53.85 7.70 54.55 11.00 ;
        RECT  56.55 7.70 57.25 11.00 ;
        RECT  0.00 11.00 60.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 4.25 ;
        RECT  1.95 2.00 2.65 3.80 ;
        RECT  4.65 2.00 5.35 3.80 ;
        RECT  7.35 2.00 8.05 3.80 ;
        RECT  10.05 2.00 10.75 3.80 ;
        RECT  12.75 2.00 13.45 3.80 ;
        RECT  15.45 2.00 16.15 3.80 ;
        RECT  18.15 2.00 18.85 3.80 ;
        RECT  20.85 2.00 21.55 3.80 ;
        RECT  58.10 2.00 59.70 4.25 ;
        RECT  0.00 0.00 60.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.30 2.45 4.00 4.80 ;
        RECT  3.45 6.75 4.15 10.55 ;
        RECT  6.00 2.45 6.70 4.80 ;
        RECT  6.15 6.75 6.85 10.55 ;
        RECT  3.45 6.75 9.55 7.25 ;
        RECT  8.70 2.45 9.40 4.80 ;
        RECT  8.85 6.75 9.55 10.55 ;
        RECT  10.20 6.75 10.90 9.60 ;
        RECT  11.40 2.45 12.10 4.80 ;
        RECT  11.55 7.70 12.25 10.55 ;
        RECT  12.90 6.75 13.60 9.60 ;
        RECT  14.10 2.45 14.80 4.80 ;
        RECT  14.25 7.70 14.95 10.55 ;
        RECT  8.85 10.05 14.95 10.55 ;
        RECT  10.20 6.75 16.30 7.25 ;
        RECT  15.60 6.75 16.30 10.55 ;
        RECT  16.80 2.45 17.50 4.80 ;
        RECT  18.30 7.70 19.00 10.55 ;
        RECT  19.50 2.45 20.20 4.80 ;
        RECT  21.00 7.70 21.70 10.55 ;
        RECT  15.60 10.05 21.70 10.55 ;
        RECT  22.20 2.45 22.90 4.80 ;
        RECT  3.30 4.30 22.90 4.80 ;
        RECT  23.55 3.40 24.25 4.10 ;
        RECT  24.90 2.45 25.60 3.15 ;
        RECT  26.25 3.40 26.95 4.10 ;
        RECT  26.70 7.70 27.40 10.55 ;
        RECT  27.60 2.45 28.30 3.15 ;
        RECT  28.95 3.40 29.65 4.10 ;
        RECT  29.40 7.70 30.10 10.55 ;
        RECT  30.30 2.45 31.00 3.15 ;
        RECT  26.70 7.70 32.80 8.20 ;
        RECT  31.65 3.40 32.35 4.10 ;
        RECT  32.10 7.70 32.80 10.55 ;
        RECT  33.00 2.45 33.70 3.15 ;
        RECT  33.45 6.75 34.15 9.60 ;
        RECT  34.35 3.40 35.05 4.10 ;
        RECT  34.80 7.70 35.50 10.55 ;
        RECT  35.70 2.45 36.40 3.15 ;
        RECT  36.15 6.75 36.85 9.60 ;
        RECT  37.05 3.40 37.75 4.10 ;
        RECT  37.50 7.70 38.20 10.55 ;
        RECT  32.10 10.05 38.20 10.55 ;
        RECT  33.45 6.75 39.35 7.25 ;
        RECT  38.40 2.45 39.10 3.15 ;
        RECT  38.85 6.75 39.35 10.55 ;
        RECT  38.85 7.70 39.55 10.55 ;
        RECT  39.75 3.40 40.45 4.10 ;
        RECT  22.20 2.45 41.80 2.95 ;
        RECT  41.10 2.45 41.80 3.15 ;
        RECT  41.55 7.70 42.25 10.55 ;
        RECT  42.45 2.45 43.15 4.10 ;
        RECT  23.55 3.60 43.15 4.10 ;
        RECT  44.25 7.70 44.95 10.55 ;
        RECT  38.85 10.05 44.95 10.55 ;
        RECT  45.15 2.45 45.85 3.15 ;
        RECT  47.10 7.70 47.80 10.55 ;
        RECT  47.85 2.45 48.55 3.15 ;
        RECT  49.80 7.70 50.50 10.55 ;
        RECT  50.55 2.45 51.25 3.15 ;
        RECT  52.50 6.75 53.20 10.55 ;
        RECT  47.10 10.05 53.20 10.55 ;
        RECT  53.25 2.45 53.95 3.15 ;
        RECT  55.20 6.75 55.90 10.55 ;
        RECT  42.45 2.45 56.65 2.95 ;
        RECT  55.95 2.45 56.65 4.10 ;
        RECT  52.50 6.75 58.60 7.25 ;
        RECT  57.90 6.75 58.60 10.55 ;
    END
END ON332X4
MACRO ON333X1
    CLASS CORE ;
    FOREIGN ON333X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.30 7.15 2.00 9.65 ;
        RECT  1.65 5.40 2.60 6.30 ;
        RECT  2.10 4.45 2.60 7.85 ;
        RECT  3.20 2.80 3.90 3.50 ;
        RECT  3.40 2.80 3.90 4.95 ;
        RECT  2.10 4.45 3.90 4.95 ;
        RECT  1.30 7.15 3.90 7.85 ;
        RECT  3.40 4.00 6.90 4.50 ;
        RECT  6.20 3.80 6.90 4.50 ;
        RECT  2.10 4.45 6.90 4.50 ;
        RECT  1.30 7.15 10.90 7.65 ;
        RECT  10.20 7.15 10.90 8.75 ;
        RECT  11.25 8.25 11.95 10.45 ;
        RECT  12.30 7.15 13.00 8.75 ;
        RECT  10.20 8.25 13.00 8.75 ;
        END
    END Q
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END J
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.25 5.35 6.30 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.25 6.80 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.35 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.25 9.60 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.20 6.35 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.75 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  13.95 5.40 15.15 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.13 ;
        PORT
        LAYER M1M ;
        RECT  15.60 5.40 16.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  6.85 8.55 7.55 11.00 ;
        RECT  15.65 7.80 16.35 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 2.05 3.80 ;
        RECT  12.95 2.00 13.65 3.30 ;
        RECT  15.65 2.00 16.35 4.45 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  8.90 3.95 15.00 4.25 ;
        RECT  4.85 2.80 5.55 3.50 ;
        RECT  7.55 2.55 8.25 3.30 ;
        RECT  4.85 2.80 8.25 3.30 ;
        RECT  8.90 3.55 9.60 4.25 ;
        RECT  7.55 2.55 10.95 3.05 ;
        RECT  4.85 2.80 10.95 3.05 ;
        RECT  10.25 2.55 10.95 3.25 ;
        RECT  11.60 2.55 12.30 4.45 ;
        RECT  8.90 3.75 12.30 4.25 ;
        RECT  14.30 2.55 15.00 4.45 ;
        RECT  11.60 3.95 15.00 4.45 ;
    END
END ON333X1
MACRO ON333X2
    CLASS CORE ;
    FOREIGN ON333X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 35.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  1.15 2.45 1.85 4.50 ;
        RECT  1.35 8.05 2.05 10.55 ;
        RECT  8.45 7.15 9.15 8.80 ;
        RECT  1.35 8.05 9.15 8.80 ;
        RECT  10.05 3.80 10.55 7.65 ;
        RECT  10.05 5.40 10.95 6.30 ;
        RECT  1.15 3.80 11.35 4.50 ;
        RECT  8.45 7.15 15.85 7.65 ;
        RECT  15.35 7.15 15.85 8.80 ;
        RECT  22.25 8.05 22.95 10.55 ;
        RECT  29.35 7.15 30.05 8.80 ;
        RECT  15.35 8.05 30.05 8.80 ;
        END
    END Q
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  4.30 5.40 5.35 6.30 ;
        END
    END J
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  5.80 5.25 6.75 6.30 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  11.40 5.40 12.35 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  21.25 5.40 22.15 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.25 20.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.25 13.75 6.35 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.30 ;
        PORT
        LAYER M1M ;
        RECT  28.25 5.40 29.25 6.35 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.28 ;
        PORT
        LAYER M1M ;
        RECT  31.05 5.35 31.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 6.28 ;
        PORT
        LAYER M1M ;
        RECT  32.40 5.40 33.35 6.35 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.35 6.55 0.85 11.00 ;
        RECT  0.35 6.55 3.45 7.25 ;
        RECT  11.80 8.10 12.50 11.00 ;
        RECT  32.70 7.10 33.40 11.00 ;
        RECT  0.00 11.00 35.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  26.00 2.00 26.70 3.55 ;
        RECT  28.70 2.00 29.40 3.55 ;
        RECT  28.70 2.85 31.85 3.55 ;
        RECT  33.85 2.00 34.55 4.45 ;
        RECT  0.00 0.00 35.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  12.00 2.45 12.70 4.50 ;
        RECT  13.50 2.45 14.20 4.50 ;
        RECT  2.50 2.45 23.70 3.15 ;
        RECT  24.35 2.45 25.05 4.50 ;
        RECT  14.85 3.80 25.05 4.50 ;
        RECT  27.35 2.45 28.05 4.50 ;
        RECT  32.50 2.55 33.20 4.50 ;
        RECT  14.85 4.00 33.20 4.50 ;
    END
END ON333X2
MACRO ON333X4
    CLASS CORE ;
    FOREIGN ON333X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 71.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  16.85 6.75 17.55 9.60 ;
        RECT  19.55 6.75 20.25 9.60 ;
        RECT  22.25 6.75 22.95 10.55 ;
        RECT  32.40 5.80 32.90 7.25 ;
        RECT  16.85 6.75 32.90 7.25 ;
        RECT  32.40 5.80 40.60 6.30 ;
        RECT  40.10 5.80 40.60 9.60 ;
        RECT  40.10 6.75 40.80 9.60 ;
        RECT  42.80 6.75 43.50 9.60 ;
        RECT  45.50 6.75 46.20 10.55 ;
        RECT  45.60 3.40 46.30 4.10 ;
        RECT  46.70 3.60 47.20 7.25 ;
        RECT  46.45 5.40 47.35 7.25 ;
        RECT  48.30 3.40 49.00 4.10 ;
        RECT  48.50 6.75 49.20 10.55 ;
        RECT  51.00 3.40 51.70 4.10 ;
        RECT  51.20 6.75 51.90 9.60 ;
        RECT  40.10 6.75 54.60 7.25 ;
        RECT  53.70 3.40 54.40 4.10 ;
        RECT  53.90 6.75 54.60 9.60 ;
        RECT  56.40 3.40 57.10 4.10 ;
        RECT  59.10 3.40 59.80 4.10 ;
        RECT  61.80 3.40 62.50 4.10 ;
        RECT  64.50 2.45 65.20 4.10 ;
        RECT  45.60 3.60 65.20 4.10 ;
        END
    END Q
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  49.25 5.40 50.15 6.30 ;
        END
    END J
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  56.25 5.40 57.15 6.30 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  63.25 5.40 64.15 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  42.25 5.40 43.15 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  31.05 5.40 31.95 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  26.85 5.40 27.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 12.60 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.50 9.55 1.20 11.00 ;
        RECT  2.00 7.15 2.70 11.00 ;
        RECT  4.70 7.70 5.40 11.00 ;
        RECT  7.40 7.70 8.10 11.00 ;
        RECT  23.75 7.70 24.45 11.00 ;
        RECT  25.25 7.70 25.95 11.00 ;
        RECT  27.95 8.65 28.65 11.00 ;
        RECT  30.65 8.70 31.35 11.00 ;
        RECT  47.00 7.70 47.70 11.00 ;
        RECT  63.35 7.70 64.05 11.00 ;
        RECT  66.05 7.70 66.75 11.00 ;
        RECT  68.75 7.25 69.45 11.00 ;
        RECT  70.25 9.60 70.95 11.00 ;
        RECT  0.00 11.00 71.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 2.95 4.25 ;
        RECT  3.75 2.00 4.45 3.80 ;
        RECT  6.45 2.00 7.15 3.80 ;
        RECT  9.15 2.00 9.85 3.80 ;
        RECT  11.85 2.00 12.55 3.80 ;
        RECT  14.55 2.00 15.25 3.80 ;
        RECT  17.25 2.00 17.95 3.80 ;
        RECT  19.95 2.00 20.65 3.80 ;
        RECT  22.65 2.00 23.35 3.80 ;
        RECT  66.20 2.00 70.50 4.25 ;
        RECT  0.00 0.00 71.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  3.35 6.75 4.05 10.55 ;
        RECT  5.10 2.45 5.80 4.80 ;
        RECT  6.05 6.75 6.75 10.55 ;
        RECT  7.80 2.45 8.50 4.80 ;
        RECT  3.35 6.75 9.45 7.25 ;
        RECT  8.75 6.75 9.45 10.55 ;
        RECT  10.10 6.75 10.80 9.60 ;
        RECT  10.50 2.45 11.20 4.80 ;
        RECT  11.45 7.70 12.15 10.55 ;
        RECT  12.80 6.75 13.50 9.60 ;
        RECT  13.20 2.45 13.90 4.80 ;
        RECT  14.15 7.70 14.85 10.55 ;
        RECT  8.75 10.05 14.85 10.55 ;
        RECT  10.10 6.75 16.20 7.25 ;
        RECT  15.50 6.75 16.20 10.55 ;
        RECT  15.90 2.45 16.60 4.80 ;
        RECT  18.20 7.70 18.90 10.55 ;
        RECT  18.60 2.45 19.30 4.80 ;
        RECT  20.90 7.70 21.60 10.55 ;
        RECT  15.50 10.05 21.60 10.55 ;
        RECT  21.30 2.45 22.00 4.80 ;
        RECT  24.00 2.45 24.70 4.80 ;
        RECT  5.10 4.30 24.70 4.80 ;
        RECT  25.35 3.40 26.05 4.10 ;
        RECT  26.60 7.70 27.30 10.55 ;
        RECT  26.70 2.45 27.40 3.15 ;
        RECT  28.05 3.40 28.75 4.10 ;
        RECT  29.30 7.70 30.00 10.55 ;
        RECT  29.40 2.45 30.10 3.15 ;
        RECT  30.75 3.40 31.45 4.10 ;
        RECT  26.60 7.70 32.70 8.20 ;
        RECT  32.00 7.70 32.70 10.55 ;
        RECT  32.10 2.45 32.80 3.15 ;
        RECT  33.35 6.75 34.05 9.60 ;
        RECT  33.45 3.40 34.15 4.10 ;
        RECT  34.70 7.70 35.40 10.55 ;
        RECT  34.80 2.45 35.50 3.15 ;
        RECT  36.05 6.75 36.75 9.60 ;
        RECT  36.15 3.40 36.85 4.10 ;
        RECT  37.40 7.70 38.10 10.55 ;
        RECT  32.00 10.05 38.10 10.55 ;
        RECT  37.50 2.45 38.20 3.15 ;
        RECT  33.35 6.75 39.45 7.25 ;
        RECT  38.75 6.75 39.45 10.55 ;
        RECT  38.85 3.40 39.55 4.10 ;
        RECT  40.20 2.45 40.90 3.15 ;
        RECT  41.45 7.70 42.15 10.55 ;
        RECT  41.55 3.40 42.25 4.10 ;
        RECT  24.00 2.45 43.60 2.95 ;
        RECT  42.90 2.45 43.60 3.15 ;
        RECT  44.15 7.70 44.85 10.55 ;
        RECT  38.75 10.05 44.85 10.55 ;
        RECT  44.25 2.45 44.95 4.10 ;
        RECT  25.35 3.60 44.95 4.10 ;
        RECT  46.95 2.45 47.65 3.15 ;
        RECT  49.65 2.45 50.35 3.15 ;
        RECT  49.85 7.70 50.55 10.55 ;
        RECT  52.35 2.45 53.05 3.15 ;
        RECT  52.55 7.70 53.25 10.55 ;
        RECT  55.05 2.45 55.75 3.15 ;
        RECT  55.25 6.75 55.95 10.55 ;
        RECT  49.85 10.05 55.95 10.55 ;
        RECT  56.60 7.70 57.30 10.55 ;
        RECT  57.75 2.45 58.45 3.15 ;
        RECT  57.95 6.75 58.65 9.60 ;
        RECT  59.30 7.70 60.00 10.55 ;
        RECT  55.25 6.75 61.35 7.25 ;
        RECT  60.45 2.45 61.15 3.15 ;
        RECT  60.65 6.75 61.35 9.60 ;
        RECT  62.00 6.75 62.70 10.55 ;
        RECT  56.60 10.05 62.70 10.55 ;
        RECT  44.25 2.45 63.85 2.95 ;
        RECT  63.15 2.45 63.85 3.15 ;
        RECT  64.70 6.75 65.40 10.55 ;
        RECT  62.00 6.75 68.10 7.25 ;
        RECT  67.40 6.75 68.10 10.55 ;
    END
END ON333X4
MACRO ON33X1
    CLASS CORE ;
    FOREIGN ON33X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.35 6.30 ;
        RECT  4.95 4.45 5.35 10.55 ;
        RECT  4.85 4.45 5.35 7.80 ;
        RECT  4.95 7.10 5.65 10.55 ;
        RECT  6.00 3.40 6.50 4.95 ;
        RECT  4.85 4.45 6.50 4.95 ;
        RECT  6.00 3.40 6.70 4.80 ;
        RECT  3.90 7.10 6.70 7.80 ;
        RECT  6.00 4.30 9.40 4.80 ;
        RECT  8.70 2.45 9.40 4.80 ;
        RECT  4.85 4.45 9.40 4.80 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.25 8.15 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.40 9.60 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.25 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.78 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.55 7.10 1.25 11.00 ;
        RECT  9.35 7.10 10.05 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.20 4.05 ;
        RECT  3.15 2.00 3.85 3.05 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 2.75 2.50 4.00 ;
        RECT  4.50 2.45 5.20 4.00 ;
        RECT  1.80 3.50 5.20 4.00 ;
        RECT  4.50 2.45 8.05 2.95 ;
        RECT  7.35 2.45 8.05 3.45 ;
    END
END ON33X1
MACRO ON33X2
    CLASS CORE ;
    FOREIGN ON33X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 26.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  10.00 7.70 10.70 10.55 ;
        RECT  12.70 6.75 13.40 10.55 ;
        RECT  12.85 3.40 13.40 10.55 ;
        RECT  10.00 10.05 13.40 10.55 ;
        RECT  12.85 3.40 13.55 4.95 ;
        RECT  12.85 5.40 13.75 6.30 ;
        RECT  12.70 6.75 16.10 7.25 ;
        RECT  15.40 6.75 16.10 9.60 ;
        RECT  15.55 3.40 16.25 4.95 ;
        RECT  18.25 3.40 18.95 4.95 ;
        RECT  20.95 3.40 21.65 4.95 ;
        RECT  12.85 4.45 21.65 4.95 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.60 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.60 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.40 18.05 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.60 ;
        PORT
        LAYER M1M ;
        RECT  21.25 5.40 22.20 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.60 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 11.00 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.60 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 5.60 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.55 6.75 1.25 11.00 ;
        RECT  0.55 6.75 3.95 7.25 ;
        RECT  3.25 6.75 3.95 9.60 ;
        RECT  22.20 7.70 22.90 11.00 ;
        RECT  24.95 7.10 25.65 11.00 ;
        RECT  0.00 11.00 26.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.80 2.00 1.50 4.00 ;
        RECT  2.65 2.00 3.35 4.00 ;
        RECT  5.35 2.00 6.05 4.00 ;
        RECT  8.05 2.00 8.75 4.00 ;
        RECT  10.75 2.00 11.45 4.00 ;
        RECT  22.45 2.00 26.00 4.00 ;
        RECT  0.00 0.00 26.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.90 7.70 2.60 10.55 ;
        RECT  4.00 2.45 4.70 4.95 ;
        RECT  4.60 6.75 5.30 10.55 ;
        RECT  1.90 10.05 5.30 10.55 ;
        RECT  5.95 7.70 6.65 10.55 ;
        RECT  4.60 6.75 8.00 7.25 ;
        RECT  6.70 2.45 7.40 4.95 ;
        RECT  7.30 6.75 8.00 9.60 ;
        RECT  8.65 6.75 9.35 10.55 ;
        RECT  5.95 10.05 9.35 10.55 ;
        RECT  9.40 2.45 10.10 4.95 ;
        RECT  8.65 6.75 12.05 7.25 ;
        RECT  11.35 6.75 12.05 9.60 ;
        RECT  11.90 2.45 12.40 4.95 ;
        RECT  4.00 4.45 12.40 4.95 ;
        RECT  14.05 7.70 14.75 10.55 ;
        RECT  14.20 2.45 14.90 3.15 ;
        RECT  16.80 6.75 17.50 10.55 ;
        RECT  14.05 10.05 17.50 10.55 ;
        RECT  16.90 2.45 17.60 3.15 ;
        RECT  18.15 7.70 18.85 10.55 ;
        RECT  16.80 6.75 20.20 7.25 ;
        RECT  11.90 2.45 20.30 2.95 ;
        RECT  19.50 6.75 20.20 9.60 ;
        RECT  19.60 2.45 20.30 3.15 ;
        RECT  20.85 6.75 21.55 10.55 ;
        RECT  18.15 10.05 21.55 10.55 ;
        RECT  20.85 6.75 24.25 7.25 ;
        RECT  23.55 6.75 24.25 10.55 ;
    END
END ON33X2
MACRO ON33X4
    CLASS CORE ;
    FOREIGN ON33X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 43.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  15.30 6.75 16.00 9.60 ;
        RECT  18.00 6.75 18.70 9.60 ;
        RECT  20.70 6.75 21.40 10.55 ;
        RECT  23.40 6.75 24.10 9.60 ;
        RECT  15.30 6.75 26.80 7.25 ;
        RECT  24.85 3.40 25.55 4.10 ;
        RECT  25.85 3.60 26.35 7.25 ;
        RECT  26.10 3.60 26.35 9.60 ;
        RECT  25.45 5.40 26.35 7.25 ;
        RECT  26.10 6.75 26.80 9.60 ;
        RECT  27.55 3.40 28.25 4.10 ;
        RECT  30.25 3.40 30.95 4.10 ;
        RECT  32.95 3.40 33.65 4.10 ;
        RECT  35.65 3.40 36.35 4.10 ;
        RECT  38.35 3.40 39.05 4.10 ;
        RECT  24.85 3.60 39.05 4.10 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 11.20 ;
        PORT
        LAYER M1M ;
        RECT  26.85 5.40 27.75 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 11.20 ;
        PORT
        LAYER M1M ;
        RECT  29.65 5.35 30.55 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 11.20 ;
        PORT
        LAYER M1M ;
        RECT  36.65 5.35 37.55 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 11.20 ;
        PORT
        LAYER M1M ;
        RECT  18.40 5.35 19.35 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 11.20 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.35 13.75 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 11.20 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.35 6.75 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 7.15 1.15 11.00 ;
        RECT  3.15 7.70 3.85 11.00 ;
        RECT  5.85 7.70 6.55 11.00 ;
        RECT  35.55 7.70 36.25 11.00 ;
        RECT  38.25 7.70 38.95 11.00 ;
        RECT  40.95 7.15 41.65 11.00 ;
        RECT  0.00 11.00 43.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.70 2.00 5.90 3.80 ;
        RECT  8.65 2.00 9.35 3.65 ;
        RECT  11.35 2.00 12.05 3.65 ;
        RECT  14.05 2.00 14.75 3.65 ;
        RECT  16.75 2.00 17.45 3.65 ;
        RECT  19.45 2.00 20.15 3.65 ;
        RECT  22.15 2.00 22.85 3.65 ;
        RECT  41.20 2.00 42.80 4.10 ;
        RECT  0.00 0.00 43.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.80 6.75 2.50 10.55 ;
        RECT  4.50 6.75 5.20 10.55 ;
        RECT  1.80 6.75 7.90 7.25 ;
        RECT  7.20 6.75 7.90 10.55 ;
        RECT  7.30 2.45 8.00 4.60 ;
        RECT  8.55 6.75 9.25 9.60 ;
        RECT  9.90 7.70 10.60 10.55 ;
        RECT  10.00 2.45 10.70 4.60 ;
        RECT  11.25 6.75 11.95 9.60 ;
        RECT  12.60 7.70 13.30 10.55 ;
        RECT  7.20 10.05 13.30 10.55 ;
        RECT  12.70 2.45 13.40 4.60 ;
        RECT  8.55 6.75 14.65 7.25 ;
        RECT  13.95 6.75 14.65 10.55 ;
        RECT  15.40 2.45 16.10 4.60 ;
        RECT  16.65 7.70 17.35 10.55 ;
        RECT  18.10 2.45 18.80 4.60 ;
        RECT  19.35 7.70 20.05 10.55 ;
        RECT  13.95 10.05 20.05 10.55 ;
        RECT  20.80 2.45 21.50 4.60 ;
        RECT  22.05 7.70 22.75 10.55 ;
        RECT  23.50 2.45 24.20 4.60 ;
        RECT  7.30 4.10 24.20 4.60 ;
        RECT  24.75 7.70 25.45 10.55 ;
        RECT  26.20 2.45 26.90 3.15 ;
        RECT  27.45 6.75 28.15 10.55 ;
        RECT  22.05 10.05 28.15 10.55 ;
        RECT  28.80 7.70 29.50 10.55 ;
        RECT  28.90 2.45 29.60 3.15 ;
        RECT  30.15 6.75 30.85 9.60 ;
        RECT  31.50 7.70 32.20 10.55 ;
        RECT  31.60 2.45 32.30 3.15 ;
        RECT  27.45 6.75 33.55 7.25 ;
        RECT  32.85 6.75 33.55 9.60 ;
        RECT  34.20 6.75 34.90 10.55 ;
        RECT  28.80 10.05 34.90 10.55 ;
        RECT  34.30 2.45 35.00 3.15 ;
        RECT  36.90 6.75 37.60 10.55 ;
        RECT  37.00 2.45 37.70 3.15 ;
        RECT  34.20 6.75 40.30 7.25 ;
        RECT  23.50 2.45 40.40 2.95 ;
        RECT  39.60 6.75 40.30 10.55 ;
        RECT  39.70 2.45 40.40 3.15 ;
    END
END ON33X4
MACRO OR2X1
    CLASS CORE ;
    FOREIGN OR2X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.15 3.10 4.95 3.80 ;
        RECT  4.45 3.10 4.95 8.95 ;
        RECT  4.25 7.15 4.95 8.95 ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  2.55 5.40 3.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 7.15 3.50 11.00 ;
        RECT  4.45 10.10 5.15 11.00 ;
        RECT  0.00 11.00 5.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 2.00 3.50 3.80 ;
        RECT  0.00 0.00 5.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.65 5.45 1.15 10.45 ;
        RECT  0.45 7.15 1.15 10.45 ;
        RECT  1.25 2.85 2.10 3.55 ;
        RECT  1.60 2.85 2.10 5.95 ;
        RECT  0.65 5.45 2.10 5.95 ;
        RECT  1.60 4.25 4.00 4.75 ;
        RECT  3.30 4.25 4.00 4.95 ;
    END
END OR2X1
MACRO OR2X2
    CLASS CORE ;
    FOREIGN OR2X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 5.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.20 2.75 4.95 4.35 ;
        RECT  4.45 2.75 4.95 10.55 ;
        RECT  4.25 8.05 4.95 10.55 ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  2.55 6.05 3.25 7.60 ;
        RECT  2.55 6.70 3.95 7.60 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.90 8.05 3.60 11.00 ;
        RECT  0.00 11.00 5.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.10 2.00 1.80 2.15 ;
        RECT  2.85 2.00 3.55 4.35 ;
        RECT  0.00 0.00 5.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.55 7.10 1.25 10.55 ;
        RECT  1.10 2.80 2.10 3.50 ;
        RECT  1.35 2.80 2.10 4.40 ;
        RECT  1.60 2.80 2.10 7.60 ;
        RECT  0.55 7.10 2.10 7.60 ;
        RECT  1.60 4.80 4.00 5.30 ;
        RECT  3.30 4.80 4.00 5.50 ;
    END
END OR2X2
MACRO OR2X3
    CLASS CORE ;
    FOREIGN OR2X3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.20 3.45 4.95 4.15 ;
        RECT  4.45 3.45 4.95 10.55 ;
        RECT  4.25 8.05 4.95 10.55 ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  2.55 6.05 3.25 7.60 ;
        RECT  2.55 6.70 3.95 7.60 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.90 8.05 3.60 11.00 ;
        RECT  5.60 8.05 6.30 11.00 ;
        RECT  0.00 11.00 7.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.10 2.00 1.80 2.15 ;
        RECT  2.85 2.00 3.55 4.15 ;
        RECT  5.55 2.00 6.25 4.15 ;
        RECT  0.00 0.00 7.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.55 7.10 1.25 10.55 ;
        RECT  1.10 2.80 2.10 3.50 ;
        RECT  1.35 2.80 2.10 4.40 ;
        RECT  1.60 2.80 2.10 7.60 ;
        RECT  0.55 7.10 2.10 7.60 ;
        RECT  1.60 4.80 4.00 5.30 ;
        RECT  3.30 4.80 4.00 5.50 ;
    END
END OR2X3
MACRO OR2X4
    CLASS CORE ;
    FOREIGN OR2X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.20 2.75 4.95 4.35 ;
        RECT  4.45 2.75 4.95 10.55 ;
        RECT  4.25 8.05 4.95 10.55 ;
        RECT  4.45 5.40 5.35 6.30 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  2.55 6.05 3.25 7.60 ;
        RECT  2.55 6.70 3.95 7.60 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.90 8.05 3.60 11.00 ;
        RECT  5.60 7.15 6.30 11.00 ;
        RECT  0.00 11.00 7.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.10 2.00 1.80 2.15 ;
        RECT  2.85 2.00 3.55 4.35 ;
        RECT  5.55 2.00 6.25 4.35 ;
        RECT  0.00 0.00 7.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.55 7.10 1.25 10.55 ;
        RECT  1.10 2.80 2.10 3.50 ;
        RECT  1.35 2.80 2.10 4.40 ;
        RECT  1.60 2.80 2.10 7.60 ;
        RECT  0.55 7.10 2.10 7.60 ;
        RECT  1.60 4.80 4.00 5.30 ;
        RECT  3.30 4.80 4.00 5.50 ;
    END
END OR2X4
MACRO OR3X1
    CLASS CORE ;
    FOREIGN OR3X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  6.95 2.55 7.85 3.25 ;
        RECT  7.25 2.55 7.65 8.95 ;
        RECT  6.95 7.15 7.65 8.95 ;
        RECT  7.25 2.55 7.85 7.75 ;
        RECT  6.95 7.15 7.85 7.75 ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.85 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.25 3.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  5.60 7.15 6.30 11.00 ;
        RECT  3.80 10.65 6.30 11.00 ;
        RECT  7.10 10.10 7.80 11.00 ;
        RECT  0.00 11.00 8.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.90 2.00 3.60 3.25 ;
        RECT  5.60 2.00 6.30 3.25 ;
        RECT  0.00 0.00 8.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 7.15 1.15 10.45 ;
        RECT  1.55 2.55 2.25 3.25 ;
        RECT  1.75 2.55 2.25 7.85 ;
        RECT  0.45 7.15 2.95 7.85 ;
        RECT  4.25 2.55 4.95 4.25 ;
        RECT  1.75 3.75 6.75 4.25 ;
        RECT  6.05 3.75 6.75 4.45 ;
    END
END OR3X1
MACRO OR3X2
    CLASS CORE ;
    FOREIGN OR3X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 8.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  7.25 2.45 7.75 10.55 ;
        RECT  6.95 7.15 7.75 10.55 ;
        RECT  7.25 2.45 7.95 4.05 ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.70 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.25 3.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  5.60 7.15 6.30 11.00 ;
        RECT  3.80 10.50 6.30 11.00 ;
        RECT  0.00 11.00 8.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.05 2.00 3.75 3.85 ;
        RECT  0.70 2.00 5.00 2.25 ;
        RECT  5.90 2.00 6.60 3.85 ;
        RECT  0.00 0.00 8.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.70 4.30 1.15 10.45 ;
        RECT  0.45 7.15 1.15 10.45 ;
        RECT  0.70 4.30 1.20 7.85 ;
        RECT  1.70 3.20 2.40 4.80 ;
        RECT  0.45 7.15 2.95 7.85 ;
        RECT  4.40 3.20 5.10 4.80 ;
        RECT  0.70 4.30 6.80 4.80 ;
        RECT  6.10 4.30 6.80 5.10 ;
    END
END OR3X2
MACRO OR3X3
    CLASS CORE ;
    FOREIGN OR3X3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  7.25 2.95 7.75 9.75 ;
        RECT  7.25 5.40 7.80 9.75 ;
        RECT  7.10 7.25 7.80 9.75 ;
        RECT  7.25 2.95 7.95 3.65 ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.70 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.25 3.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  5.60 7.25 6.30 11.00 ;
        RECT  3.80 10.50 6.30 11.00 ;
        RECT  8.45 7.25 9.15 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.05 2.00 3.75 3.85 ;
        RECT  0.50 2.00 4.80 2.25 ;
        RECT  5.90 2.00 6.60 3.65 ;
        RECT  8.60 2.00 9.30 3.65 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.70 4.30 1.15 10.45 ;
        RECT  0.45 7.15 1.15 10.45 ;
        RECT  0.70 4.30 1.20 7.85 ;
        RECT  1.70 3.20 2.40 4.80 ;
        RECT  0.45 7.15 2.95 7.85 ;
        RECT  4.40 3.20 5.10 4.80 ;
        RECT  0.70 4.30 6.80 4.80 ;
        RECT  6.10 4.30 6.80 5.10 ;
    END
END OR3X3
MACRO OR3X4
    CLASS CORE ;
    FOREIGN OR3X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  7.25 2.45 7.75 10.55 ;
        RECT  6.95 7.15 7.75 10.55 ;
        RECT  7.25 2.45 7.95 4.05 ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.70 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.25 3.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  5.60 7.15 6.30 11.00 ;
        RECT  3.80 10.50 6.30 11.00 ;
        RECT  8.30 7.15 9.00 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.05 2.00 3.75 3.85 ;
        RECT  0.50 2.00 4.80 2.25 ;
        RECT  5.90 2.00 6.60 3.85 ;
        RECT  8.60 2.00 9.30 3.85 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.70 4.30 1.15 10.45 ;
        RECT  0.45 7.15 1.15 10.45 ;
        RECT  0.70 4.30 1.20 7.85 ;
        RECT  1.70 3.20 2.40 4.80 ;
        RECT  0.45 7.15 2.95 7.85 ;
        RECT  4.40 3.20 5.10 4.80 ;
        RECT  0.70 4.30 6.80 4.80 ;
        RECT  6.10 4.30 6.80 5.10 ;
    END
END OR3X4
MACRO OR4X1
    CLASS CORE ;
    FOREIGN OR4X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.90 3.60 5.40 8.85 ;
        RECT  4.70 7.25 5.40 8.85 ;
        RECT  5.65 2.45 6.35 4.10 ;
        RECT  4.90 3.60 6.35 4.10 ;
        RECT  5.65 2.80 6.75 3.70 ;
        RECT  4.90 3.60 6.75 3.70 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.35 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  7.25 4.10 8.15 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.30 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.20 7.70 3.90 11.00 ;
        RECT  6.20 7.45 6.90 11.00 ;
        RECT  10.05 9.55 10.75 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.75 ;
        RECT  3.30 2.00 4.00 3.90 ;
        RECT  7.35 2.00 8.05 3.65 ;
        RECT  10.05 2.00 10.75 3.65 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.85 6.75 1.55 10.55 ;
        RECT  1.80 3.05 2.50 3.75 ;
        RECT  2.00 3.05 2.50 4.85 ;
        RECT  2.00 4.35 3.65 4.85 ;
        RECT  3.15 4.35 3.65 7.25 ;
        RECT  0.85 6.75 3.65 7.25 ;
        RECT  3.15 5.25 4.45 5.95 ;
        RECT  5.85 5.25 6.55 5.95 ;
        RECT  5.85 5.45 9.25 5.95 ;
        RECT  8.75 3.00 9.25 10.55 ;
        RECT  8.55 7.15 9.25 10.55 ;
        RECT  8.70 3.00 9.40 3.70 ;
    END
END OR4X1
MACRO OR4X2
    CLASS CORE ;
    FOREIGN OR4X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 11.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  5.05 3.95 5.55 10.55 ;
        RECT  4.85 7.15 5.55 10.55 ;
        RECT  5.65 2.80 6.35 4.45 ;
        RECT  5.05 3.95 6.35 4.45 ;
        RECT  5.65 2.80 6.75 3.70 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.40 10.95 6.35 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  7.25 4.10 8.15 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.25 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.50 7.70 4.20 11.00 ;
        RECT  6.20 7.45 6.90 11.00 ;
        RECT  10.05 9.55 10.75 11.00 ;
        RECT  0.00 11.00 11.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.75 ;
        RECT  3.30 2.00 4.00 3.85 ;
        RECT  7.35 2.00 8.05 3.65 ;
        RECT  10.05 2.00 10.75 3.65 ;
        RECT  0.00 0.00 11.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.15 6.75 1.85 10.55 ;
        RECT  1.80 3.05 2.50 3.75 ;
        RECT  2.00 3.05 2.50 4.80 ;
        RECT  2.00 4.30 3.65 4.80 ;
        RECT  3.15 4.30 3.65 7.25 ;
        RECT  1.15 6.75 3.65 7.25 ;
        RECT  3.15 5.25 4.60 5.95 ;
        RECT  6.00 5.25 6.70 5.95 ;
        RECT  6.00 5.45 9.25 5.95 ;
        RECT  8.75 3.00 9.25 10.55 ;
        RECT  8.55 7.15 9.25 10.55 ;
        RECT  8.70 3.00 9.40 3.70 ;
    END
END OR4X2
MACRO OR4X3
    CLASS CORE ;
    FOREIGN OR4X3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.70 7.70 5.40 10.50 ;
        RECT  5.85 3.15 6.35 8.20 ;
        RECT  5.85 3.15 6.75 5.00 ;
        RECT  4.70 7.70 8.10 8.20 ;
        RECT  7.40 7.70 8.10 10.55 ;
        RECT  8.25 2.45 8.75 3.90 ;
        RECT  5.65 3.15 8.75 3.90 ;
        RECT  8.25 2.45 8.95 3.15 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.25 10.95 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.25 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.20 7.70 3.90 11.00 ;
        RECT  6.05 8.65 6.75 11.00 ;
        RECT  8.90 7.70 9.60 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.75 ;
        RECT  3.30 2.00 4.00 3.85 ;
        RECT  11.75 2.00 12.25 4.50 ;
        RECT  10.70 3.80 12.25 4.50 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.85 6.75 1.55 10.55 ;
        RECT  1.80 3.05 2.50 3.75 ;
        RECT  2.00 3.05 2.50 4.80 ;
        RECT  2.00 4.30 3.65 4.80 ;
        RECT  3.15 4.30 3.65 7.25 ;
        RECT  0.85 6.75 3.65 7.25 ;
        RECT  3.15 5.25 4.50 5.95 ;
        RECT  7.85 6.55 8.55 7.25 ;
        RECT  9.10 4.30 9.60 7.25 ;
        RECT  9.60 2.65 10.10 4.80 ;
        RECT  9.10 4.30 10.10 4.80 ;
        RECT  7.85 6.75 11.95 7.25 ;
        RECT  10.60 2.45 11.30 3.15 ;
        RECT  9.60 2.65 11.30 3.15 ;
        RECT  11.25 6.75 11.95 10.55 ;
    END
END OR4X3
MACRO OR4X4
    CLASS CORE ;
    FOREIGN OR4X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.15 6.50 4.85 10.55 ;
        RECT  5.85 3.20 6.75 5.00 ;
        RECT  6.25 3.20 6.75 7.00 ;
        RECT  4.15 6.50 7.55 7.00 ;
        RECT  6.85 6.50 7.55 10.55 ;
        RECT  5.65 3.20 10.55 3.90 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  11.45 4.10 12.35 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.35 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.25 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 7.70 3.50 11.00 ;
        RECT  5.50 7.45 6.20 11.00 ;
        RECT  8.20 7.45 8.90 11.00 ;
        RECT  10.05 7.40 10.75 11.00 ;
        RECT  14.25 7.45 14.95 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.75 ;
        RECT  3.30 2.00 4.00 3.85 ;
        RECT  11.55 2.00 12.25 3.65 ;
        RECT  14.25 2.00 14.95 3.65 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 6.75 1.15 10.55 ;
        RECT  1.80 3.05 2.50 3.75 ;
        RECT  2.00 3.05 2.50 4.80 ;
        RECT  2.00 4.30 3.65 4.80 ;
        RECT  3.15 4.30 3.65 7.25 ;
        RECT  0.45 6.75 3.65 7.25 ;
        RECT  3.15 4.80 4.45 5.50 ;
        RECT  8.00 5.25 8.70 5.95 ;
        RECT  12.10 5.45 12.60 10.55 ;
        RECT  11.90 7.15 12.60 10.55 ;
        RECT  12.95 3.00 13.45 5.95 ;
        RECT  8.00 5.45 13.45 5.95 ;
        RECT  12.90 3.00 13.60 3.70 ;
    END
END OR4X4
MACRO OR5X1
    CLASS CORE ;
    FOREIGN OR5X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  7.15 2.45 7.45 9.25 ;
        RECT  6.75 7.55 7.45 9.25 ;
        RECT  7.15 2.45 7.65 8.05 ;
        RECT  6.75 7.55 7.65 8.05 ;
        RECT  7.15 2.45 7.85 4.15 ;
        RECT  7.15 2.80 8.15 3.70 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.40 9.55 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.43 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.45 5.35 7.60 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  5.25 8.10 5.95 11.00 ;
        RECT  6.75 10.30 7.45 11.00 ;
        RECT  8.25 7.35 8.95 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.95 2.00 2.65 4.00 ;
        RECT  4.80 2.00 5.50 4.00 ;
        RECT  8.75 2.00 9.45 3.75 ;
        RECT  11.45 2.00 12.15 3.75 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  10.50 3.05 10.80 7.70 ;
        RECT  10.50 7.15 11.30 7.70 ;
        RECT  0.45 7.55 1.15 10.45 ;
        RECT  0.60 3.30 1.30 4.95 ;
        RECT  2.05 4.45 2.55 8.25 ;
        RECT  0.45 7.55 2.55 8.25 ;
        RECT  3.30 3.30 4.00 4.95 ;
        RECT  0.60 4.45 6.15 4.95 ;
        RECT  5.45 4.45 6.15 5.35 ;
        RECT  8.30 4.20 9.00 4.90 ;
        RECT  8.30 4.20 11.00 4.70 ;
        RECT  10.60 3.05 10.80 10.55 ;
        RECT  10.10 3.05 10.80 4.70 ;
        RECT  10.60 4.20 11.00 10.55 ;
        RECT  10.50 4.20 11.00 7.70 ;
        RECT  10.60 7.15 11.30 10.55 ;
    END
END OR5X1
MACRO OR5X2
    CLASS CORE ;
    FOREIGN OR5X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  6.55 4.00 7.05 10.55 ;
        RECT  6.55 7.15 7.25 10.55 ;
        RECT  7.15 2.80 7.85 4.50 ;
        RECT  6.55 4.00 7.85 4.50 ;
        RECT  7.15 2.80 8.15 3.70 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  11.45 5.40 12.35 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.55 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.35 3.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.20 5.35 7.60 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  5.15 8.10 5.85 11.00 ;
        RECT  7.90 7.35 8.60 11.00 ;
        RECT  0.00 11.00 12.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.90 2.00 2.60 3.95 ;
        RECT  4.75 2.00 5.45 3.95 ;
        RECT  8.75 2.00 9.45 3.65 ;
        RECT  11.45 2.00 12.15 3.65 ;
        RECT  0.00 0.00 12.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 7.55 1.15 10.45 ;
        RECT  0.55 3.35 1.25 4.90 ;
        RECT  1.95 4.40 2.45 8.25 ;
        RECT  0.45 7.55 2.45 8.25 ;
        RECT  3.25 3.35 3.95 4.90 ;
        RECT  0.55 4.40 6.00 4.90 ;
        RECT  5.30 4.40 6.00 5.55 ;
        RECT  7.50 5.70 8.20 6.40 ;
        RECT  10.10 3.00 10.95 3.70 ;
        RECT  7.50 5.70 10.95 6.20 ;
        RECT  10.45 3.00 10.95 10.55 ;
        RECT  10.25 7.15 10.95 10.55 ;
    END
END OR5X2
MACRO OR5X3
    CLASS CORE ;
    FOREIGN OR5X3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  6.65 6.60 7.35 9.80 ;
        RECT  7.25 3.15 8.15 5.00 ;
        RECT  7.65 3.15 8.15 7.10 ;
        RECT  6.65 6.60 10.05 7.10 ;
        RECT  9.35 6.60 10.05 9.80 ;
        RECT  10.05 2.45 10.75 3.90 ;
        RECT  7.25 3.15 10.75 3.90 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  11.45 4.10 12.35 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.20 5.35 7.60 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  5.15 8.10 5.85 11.00 ;
        RECT  8.00 7.55 8.70 11.00 ;
        RECT  10.85 7.55 11.55 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.25 2.00 2.95 4.00 ;
        RECT  5.10 2.00 5.80 4.00 ;
        RECT  11.55 2.00 12.25 3.65 ;
        RECT  14.25 2.00 14.95 3.65 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.90 3.35 1.15 10.45 ;
        RECT  0.45 7.25 1.15 10.45 ;
        RECT  0.90 3.35 1.20 7.95 ;
        RECT  0.70 4.45 1.20 7.95 ;
        RECT  0.90 3.35 1.60 4.95 ;
        RECT  0.45 7.25 2.45 7.95 ;
        RECT  3.60 3.35 4.30 4.95 ;
        RECT  0.70 4.45 6.10 4.95 ;
        RECT  5.40 4.45 6.10 5.55 ;
        RECT  9.80 5.45 10.50 6.15 ;
        RECT  12.90 3.00 13.70 3.70 ;
        RECT  9.80 5.45 13.70 5.95 ;
        RECT  13.20 3.00 13.70 10.55 ;
        RECT  13.20 7.15 13.90 10.55 ;
    END
END OR5X3
MACRO OR5X4
    CLASS CORE ;
    FOREIGN OR5X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  6.50 6.50 7.20 10.55 ;
        RECT  7.25 3.20 8.15 5.00 ;
        RECT  7.65 3.20 8.15 7.00 ;
        RECT  6.50 6.50 9.90 7.00 ;
        RECT  9.20 6.50 9.90 10.55 ;
        RECT  7.25 3.20 12.15 3.90 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  12.85 4.10 13.75 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.05 5.35 7.60 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  5.15 8.10 5.85 11.00 ;
        RECT  7.85 7.45 8.55 11.00 ;
        RECT  10.55 7.45 11.25 11.00 ;
        RECT  15.65 7.45 16.35 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.05 2.00 2.75 4.00 ;
        RECT  4.90 2.00 5.60 4.00 ;
        RECT  12.95 2.00 13.65 3.65 ;
        RECT  15.65 2.00 16.35 3.65 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.70 3.35 1.15 10.45 ;
        RECT  0.45 7.25 1.15 10.45 ;
        RECT  0.70 3.35 1.20 7.95 ;
        RECT  0.70 3.35 1.40 4.95 ;
        RECT  0.45 7.25 2.45 7.95 ;
        RECT  3.40 3.35 4.10 4.95 ;
        RECT  0.70 4.45 6.25 4.95 ;
        RECT  5.55 4.45 6.25 5.50 ;
        RECT  9.65 5.25 10.35 5.95 ;
        RECT  13.50 5.45 14.00 10.55 ;
        RECT  13.30 7.15 14.00 10.55 ;
        RECT  14.30 3.00 14.80 5.95 ;
        RECT  9.65 5.45 14.80 5.95 ;
        RECT  14.30 3.00 15.00 3.70 ;
    END
END OR5X4
MACRO OR6X1
    CLASS CORE ;
    FOREIGN OR6X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 15.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.45 6.70 5.00 10.25 ;
        RECT  4.85 3.55 5.00 10.25 ;
        RECT  4.30 8.65 5.00 10.25 ;
        RECT  4.85 3.55 5.35 8.20 ;
        RECT  4.45 6.70 5.35 8.20 ;
        RECT  4.45 7.70 7.70 8.20 ;
        RECT  6.65 2.45 7.35 4.05 ;
        RECT  4.85 3.55 7.35 4.05 ;
        RECT  7.00 7.70 7.70 10.20 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  10.05 5.25 10.95 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  8.65 5.40 9.55 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.25 13.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.40 15.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.30 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 7.70 3.50 11.00 ;
        RECT  5.65 8.65 6.35 11.00 ;
        RECT  11.80 8.30 12.50 11.00 ;
        RECT  0.00 11.00 15.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.15 ;
        RECT  3.30 2.00 4.00 3.90 ;
        RECT  8.85 2.00 9.55 3.75 ;
        RECT  11.55 2.00 12.25 3.75 ;
        RECT  14.25 2.00 14.95 3.80 ;
        RECT  0.00 0.00 15.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 6.75 1.15 10.55 ;
        RECT  1.80 2.45 2.50 3.15 ;
        RECT  2.00 2.45 2.50 4.85 ;
        RECT  2.00 4.35 3.50 4.85 ;
        RECT  3.00 4.35 3.50 7.25 ;
        RECT  0.45 6.75 3.50 7.25 ;
        RECT  3.00 4.85 4.30 5.55 ;
        RECT  6.20 4.50 6.90 5.25 ;
        RECT  6.20 4.50 8.20 5.00 ;
        RECT  7.70 4.45 8.20 7.25 ;
        RECT  8.15 9.85 8.85 10.55 ;
        RECT  8.60 4.30 9.10 4.95 ;
        RECT  6.20 4.50 9.10 4.95 ;
        RECT  7.70 6.75 10.15 7.25 ;
        RECT  9.45 6.75 10.15 9.60 ;
        RECT  8.60 4.30 10.70 4.80 ;
        RECT  7.70 4.45 10.70 4.80 ;
        RECT  10.20 3.05 10.70 4.80 ;
        RECT  6.20 4.50 10.70 4.80 ;
        RECT  10.20 3.05 10.90 3.75 ;
        RECT  10.75 7.15 11.25 10.55 ;
        RECT  8.15 10.05 11.25 10.55 ;
        RECT  11.80 4.30 12.30 7.65 ;
        RECT  12.90 3.05 13.40 4.80 ;
        RECT  11.80 4.30 13.40 4.80 ;
        RECT  12.90 3.05 13.60 3.75 ;
        RECT  10.75 7.15 14.85 7.65 ;
        RECT  14.15 7.15 14.85 10.55 ;
    END
END OR6X1
MACRO OR6X2
    CLASS CORE ;
    FOREIGN OR6X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.30 7.70 5.00 10.15 ;
        RECT  7.65 4.45 7.70 10.15 ;
        RECT  7.00 7.70 7.70 10.15 ;
        RECT  7.65 4.45 8.15 8.20 ;
        RECT  7.25 6.70 8.15 8.20 ;
        RECT  4.30 7.70 10.40 8.20 ;
        RECT  9.70 7.70 10.40 10.15 ;
        RECT  8.70 4.25 11.45 4.95 ;
        RECT  10.75 2.45 11.45 4.95 ;
        RECT  7.65 4.45 11.45 4.95 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.25 15.15 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.25 17.95 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.40 19.35 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.30 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 7.70 3.50 11.00 ;
        RECT  5.65 8.65 6.35 11.00 ;
        RECT  8.35 8.65 9.05 11.00 ;
        RECT  11.05 8.65 11.75 11.00 ;
        RECT  16.00 8.30 16.70 11.00 ;
        RECT  0.00 11.00 19.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.65 ;
        RECT  3.15 2.00 3.85 3.65 ;
        RECT  5.35 2.00 6.05 4.25 ;
        RECT  13.05 2.00 13.75 3.75 ;
        RECT  15.75 2.00 16.45 3.75 ;
        RECT  18.45 2.00 19.15 3.80 ;
        RECT  0.00 0.00 19.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 6.75 1.15 10.55 ;
        RECT  1.80 2.95 2.50 3.65 ;
        RECT  2.00 2.95 2.50 4.70 ;
        RECT  2.00 4.20 3.50 4.70 ;
        RECT  3.00 4.20 3.50 7.25 ;
        RECT  0.45 6.75 3.50 7.25 ;
        RECT  3.00 6.25 5.90 6.75 ;
        RECT  5.20 6.05 5.90 6.75 ;
        RECT  9.25 6.55 9.95 7.25 ;
        RECT  9.25 6.55 12.40 7.05 ;
        RECT  11.90 4.30 12.40 7.60 ;
        RECT  12.20 9.85 12.90 10.55 ;
        RECT  11.90 7.10 14.35 7.60 ;
        RECT  13.65 7.10 14.35 9.60 ;
        RECT  14.40 3.05 14.90 4.80 ;
        RECT  11.90 4.30 14.90 4.80 ;
        RECT  14.40 3.05 15.10 3.75 ;
        RECT  14.95 7.15 15.45 10.55 ;
        RECT  12.20 10.05 15.45 10.55 ;
        RECT  16.00 4.30 16.50 7.65 ;
        RECT  17.10 3.05 17.60 4.80 ;
        RECT  16.00 4.30 17.60 4.80 ;
        RECT  17.10 3.05 17.80 3.75 ;
        RECT  14.95 7.15 19.05 7.65 ;
        RECT  18.35 7.15 19.05 10.55 ;
    END
END OR6X2
MACRO OR6X3
    CLASS CORE ;
    FOREIGN OR6X3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.30 7.40 5.00 10.55 ;
        RECT  7.25 4.10 8.15 5.00 ;
        RECT  7.65 4.10 7.70 10.55 ;
        RECT  7.00 7.40 7.70 10.55 ;
        RECT  7.65 4.10 8.15 7.90 ;
        RECT  4.30 7.40 10.40 7.90 ;
        RECT  9.70 7.40 10.40 10.55 ;
        RECT  10.95 2.45 11.45 4.80 ;
        RECT  6.65 4.10 11.45 4.80 ;
        RECT  10.95 2.45 12.25 3.15 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.25 15.15 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.25 17.95 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.40 19.35 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.30 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 7.90 3.50 11.00 ;
        RECT  5.65 8.35 6.35 11.00 ;
        RECT  8.35 8.35 9.05 11.00 ;
        RECT  11.05 8.35 11.75 11.00 ;
        RECT  16.00 8.30 16.70 11.00 ;
        RECT  0.00 11.00 19.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.65 ;
        RECT  3.30 2.00 4.00 3.70 ;
        RECT  13.05 2.00 13.75 3.75 ;
        RECT  15.75 2.00 16.45 3.75 ;
        RECT  18.45 2.00 19.15 3.80 ;
        RECT  0.00 0.00 19.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 6.75 1.15 10.55 ;
        RECT  1.80 2.95 2.50 3.65 ;
        RECT  2.00 2.95 2.50 4.85 ;
        RECT  2.00 4.35 3.50 4.85 ;
        RECT  3.00 4.35 3.50 7.25 ;
        RECT  0.45 6.75 3.50 7.25 ;
        RECT  3.00 6.25 4.45 6.95 ;
        RECT  0.45 6.75 4.45 6.95 ;
        RECT  10.15 5.80 10.85 6.50 ;
        RECT  10.15 5.80 12.40 6.30 ;
        RECT  11.90 4.30 12.40 7.60 ;
        RECT  12.20 9.85 12.90 10.55 ;
        RECT  11.90 7.10 14.35 7.60 ;
        RECT  13.65 7.10 14.35 9.60 ;
        RECT  14.40 3.05 14.90 4.80 ;
        RECT  11.90 4.30 14.90 4.80 ;
        RECT  14.40 3.05 15.10 3.75 ;
        RECT  14.95 7.15 15.45 10.55 ;
        RECT  12.20 10.05 15.45 10.55 ;
        RECT  16.00 4.30 16.50 7.65 ;
        RECT  17.10 3.05 17.60 4.80 ;
        RECT  16.00 4.30 17.60 4.80 ;
        RECT  17.10 3.05 17.80 3.75 ;
        RECT  14.95 7.15 19.05 7.65 ;
        RECT  18.35 7.15 19.05 10.55 ;
    END
END OR6X3
MACRO OR6X4
    CLASS CORE ;
    FOREIGN OR6X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.50 7.60 5.00 10.55 ;
        RECT  4.30 8.90 5.00 10.55 ;
        RECT  6.50 4.10 7.00 8.10 ;
        RECT  7.00 7.60 7.50 10.55 ;
        RECT  7.00 8.90 7.70 10.55 ;
        RECT  6.50 4.10 8.15 5.00 ;
        RECT  4.50 7.60 10.20 8.10 ;
        RECT  9.70 7.60 10.20 10.55 ;
        RECT  9.70 8.95 10.40 10.55 ;
        RECT  13.75 2.45 14.25 4.80 ;
        RECT  6.50 4.10 14.25 4.80 ;
        RECT  13.75 2.45 15.05 3.15 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.25 17.95 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.25 20.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  21.25 5.40 22.15 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.30 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 8.30 3.50 11.00 ;
        RECT  5.65 8.55 6.35 11.00 ;
        RECT  8.35 8.55 9.05 11.00 ;
        RECT  11.05 8.35 11.75 11.00 ;
        RECT  12.55 9.20 15.05 11.00 ;
        RECT  18.80 8.30 19.50 11.00 ;
        RECT  0.00 11.00 22.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.65 ;
        RECT  3.30 2.00 4.00 3.70 ;
        RECT  15.85 2.00 16.55 3.75 ;
        RECT  18.55 2.00 19.25 3.75 ;
        RECT  21.25 2.00 21.95 3.80 ;
        RECT  0.00 0.00 22.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.65 6.75 1.15 10.55 ;
        RECT  0.45 8.50 1.15 10.55 ;
        RECT  1.80 2.95 2.50 3.65 ;
        RECT  2.00 2.95 2.50 4.85 ;
        RECT  2.00 4.35 3.50 4.85 ;
        RECT  3.00 4.35 3.50 7.25 ;
        RECT  0.65 6.75 3.50 7.25 ;
        RECT  3.00 6.25 4.45 6.95 ;
        RECT  0.65 6.75 4.45 6.95 ;
        RECT  7.45 6.45 8.15 7.15 ;
        RECT  10.15 5.50 10.85 6.20 ;
        RECT  7.45 6.65 14.25 7.15 ;
        RECT  13.75 6.65 14.25 8.65 ;
        RECT  10.15 5.50 15.20 6.00 ;
        RECT  14.70 4.30 15.20 7.60 ;
        RECT  13.75 8.15 16.00 8.65 ;
        RECT  15.50 8.15 16.00 10.55 ;
        RECT  14.70 7.10 17.15 7.60 ;
        RECT  16.45 7.10 17.15 9.60 ;
        RECT  17.20 3.05 17.70 4.80 ;
        RECT  14.70 4.30 17.70 4.80 ;
        RECT  17.20 3.05 17.90 3.75 ;
        RECT  17.75 7.15 18.25 10.55 ;
        RECT  15.50 10.05 18.25 10.55 ;
        RECT  18.80 4.30 19.30 7.65 ;
        RECT  19.90 3.05 20.40 4.80 ;
        RECT  18.80 4.30 20.40 4.80 ;
        RECT  19.90 3.05 20.60 3.75 ;
        RECT  17.75 7.15 21.85 7.65 ;
        RECT  21.15 7.15 21.85 10.55 ;
    END
END OR6X4
MACRO OR7X1
    CLASS CORE ;
    FOREIGN OR7X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.45 4.10 5.35 5.00 ;
        RECT  4.15 7.70 4.85 10.15 ;
        RECT  4.85 4.10 5.35 8.20 ;
        RECT  4.15 7.70 7.55 8.20 ;
        RECT  6.50 2.45 7.20 4.60 ;
        RECT  4.45 4.10 7.20 4.60 ;
        RECT  6.85 7.70 7.55 10.15 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.25 15.15 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  11.45 4.10 12.35 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  10.05 4.10 10.95 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  8.65 4.10 9.55 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.30 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 8.55 3.50 11.00 ;
        RECT  5.50 8.65 6.20 11.00 ;
        RECT  13.20 8.20 13.90 11.00 ;
        RECT  0.00 11.00 16.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.65 ;
        RECT  3.15 2.00 3.85 3.60 ;
        RECT  10.10 2.00 10.80 2.70 ;
        RECT  12.95 2.00 13.65 3.10 ;
        RECT  15.65 2.00 16.35 3.15 ;
        RECT  0.00 0.00 16.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 6.75 1.15 10.55 ;
        RECT  1.80 2.95 2.50 3.65 ;
        RECT  2.00 2.95 2.50 4.70 ;
        RECT  2.00 4.20 3.50 4.70 ;
        RECT  3.00 4.20 3.50 7.25 ;
        RECT  0.45 6.75 3.50 7.25 ;
        RECT  3.00 6.05 4.40 6.75 ;
        RECT  5.80 5.60 6.50 6.30 ;
        RECT  7.20 6.55 8.50 7.25 ;
        RECT  7.70 3.15 8.20 6.10 ;
        RECT  8.00 6.55 8.50 10.55 ;
        RECT  8.60 2.45 9.30 3.65 ;
        RECT  5.80 5.60 10.35 6.10 ;
        RECT  9.85 5.60 10.35 9.15 ;
        RECT  9.85 7.10 10.55 9.15 ;
        RECT  8.95 8.45 10.55 9.15 ;
        RECT  11.60 2.45 12.30 3.65 ;
        RECT  7.70 3.15 12.30 3.65 ;
        RECT  12.15 7.15 12.65 10.55 ;
        RECT  8.00 10.05 12.65 10.55 ;
        RECT  13.20 4.30 13.70 7.65 ;
        RECT  14.30 2.45 14.80 4.80 ;
        RECT  13.20 4.30 14.80 4.80 ;
        RECT  14.30 2.45 15.00 3.15 ;
        RECT  12.15 7.15 16.25 7.65 ;
        RECT  15.55 7.15 16.25 10.55 ;
    END
END OR7X1
MACRO OR7X2
    CLASS CORE ;
    FOREIGN OR7X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.30 7.70 5.00 10.15 ;
        RECT  6.75 4.50 7.25 8.20 ;
        RECT  7.00 7.70 7.70 10.15 ;
        RECT  7.25 4.10 8.15 5.00 ;
        RECT  4.30 7.70 10.40 8.20 ;
        RECT  9.70 7.70 10.40 10.15 ;
        RECT  7.25 4.25 11.45 5.00 ;
        RECT  10.75 2.45 11.45 5.00 ;
        RECT  6.75 4.50 11.45 5.00 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.25 19.35 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  15.65 4.10 16.55 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  14.25 4.10 15.15 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  12.85 4.10 13.75 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.30 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 7.70 3.50 11.00 ;
        RECT  5.65 8.65 6.35 11.00 ;
        RECT  8.35 8.65 9.05 11.00 ;
        RECT  11.05 8.65 11.75 11.00 ;
        RECT  17.25 8.20 17.95 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.65 ;
        RECT  3.15 2.00 3.85 3.65 ;
        RECT  5.35 2.00 6.05 4.25 ;
        RECT  14.30 2.00 15.00 2.70 ;
        RECT  17.15 2.00 17.85 3.10 ;
        RECT  19.85 2.00 20.55 3.15 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 6.75 1.15 10.55 ;
        RECT  1.80 2.95 2.50 3.65 ;
        RECT  2.00 2.95 2.50 4.70 ;
        RECT  2.00 4.20 3.50 4.70 ;
        RECT  3.00 4.20 3.50 7.25 ;
        RECT  0.45 6.75 3.50 7.25 ;
        RECT  3.00 6.25 5.90 6.75 ;
        RECT  5.20 6.05 5.90 6.75 ;
        RECT  7.70 6.55 8.40 7.25 ;
        RECT  11.90 3.15 12.40 7.05 ;
        RECT  12.20 9.85 12.90 10.55 ;
        RECT  12.80 2.45 13.50 3.65 ;
        RECT  7.70 6.55 14.40 7.05 ;
        RECT  13.90 6.55 14.40 9.15 ;
        RECT  13.90 7.10 14.60 9.15 ;
        RECT  13.00 8.45 14.60 9.15 ;
        RECT  15.80 2.45 16.50 3.65 ;
        RECT  11.90 3.15 16.50 3.65 ;
        RECT  16.20 7.15 16.70 10.55 ;
        RECT  12.20 10.05 16.70 10.55 ;
        RECT  17.40 4.30 17.90 7.65 ;
        RECT  18.50 2.45 19.00 4.80 ;
        RECT  17.40 4.30 19.00 4.80 ;
        RECT  18.50 2.45 19.20 3.15 ;
        RECT  16.20 7.15 20.45 7.65 ;
        RECT  19.75 7.15 20.45 10.55 ;
    END
END OR7X2
MACRO OR7X3
    CLASS CORE ;
    FOREIGN OR7X3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.30 7.40 5.00 10.55 ;
        RECT  7.05 4.10 7.55 10.55 ;
        RECT  7.00 7.40 7.70 10.55 ;
        RECT  7.05 4.10 8.15 5.00 ;
        RECT  4.30 7.40 10.40 7.90 ;
        RECT  9.70 7.40 10.40 10.55 ;
        RECT  10.95 2.45 11.45 4.80 ;
        RECT  6.65 4.10 11.45 4.80 ;
        RECT  10.95 2.45 12.25 3.15 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.25 19.35 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.40 20.75 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  16.35 4.45 16.85 6.30 ;
        RECT  15.65 5.40 16.85 6.30 ;
        RECT  16.35 4.45 17.05 5.15 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  14.25 5.10 15.15 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  12.85 5.40 13.75 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.30 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 7.90 3.50 11.00 ;
        RECT  5.65 8.35 6.35 11.00 ;
        RECT  8.35 8.35 9.05 11.00 ;
        RECT  11.05 8.35 11.75 11.00 ;
        RECT  17.25 8.20 17.95 11.00 ;
        RECT  0.00 11.00 21.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.65 ;
        RECT  3.30 2.00 4.00 3.70 ;
        RECT  14.45 2.00 15.15 3.05 ;
        RECT  17.15 2.00 17.85 3.10 ;
        RECT  19.85 2.00 20.55 3.10 ;
        RECT  0.00 0.00 21.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 6.75 1.15 10.55 ;
        RECT  1.80 2.95 2.50 3.65 ;
        RECT  2.00 2.95 2.50 4.85 ;
        RECT  2.00 4.35 3.50 4.85 ;
        RECT  3.00 4.35 3.50 7.25 ;
        RECT  0.45 6.75 3.50 7.25 ;
        RECT  3.00 6.25 4.45 6.95 ;
        RECT  0.45 6.75 4.45 6.95 ;
        RECT  8.00 6.25 8.70 6.95 ;
        RECT  11.90 3.60 12.40 7.25 ;
        RECT  8.00 6.25 12.40 6.75 ;
        RECT  12.20 9.85 12.90 10.55 ;
        RECT  13.10 2.45 13.80 4.10 ;
        RECT  11.90 3.60 13.80 4.10 ;
        RECT  11.90 6.75 14.60 7.25 ;
        RECT  13.90 6.75 14.60 9.15 ;
        RECT  13.00 8.45 14.60 9.15 ;
        RECT  13.10 3.50 16.30 4.00 ;
        RECT  15.80 2.45 16.30 4.00 ;
        RECT  11.90 3.60 16.30 4.00 ;
        RECT  15.80 2.45 16.50 3.15 ;
        RECT  16.20 7.15 16.70 10.55 ;
        RECT  12.20 10.05 16.70 10.55 ;
        RECT  17.50 4.30 18.00 7.65 ;
        RECT  18.50 2.45 19.00 4.80 ;
        RECT  17.50 4.30 19.00 4.80 ;
        RECT  18.50 2.45 19.20 3.15 ;
        RECT  16.20 7.15 20.45 7.65 ;
        RECT  19.75 7.15 20.45 10.55 ;
    END
END OR7X3
MACRO OR7X4
    CLASS CORE ;
    FOREIGN OR7X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  4.50 7.60 5.00 10.55 ;
        RECT  4.30 8.90 5.00 10.55 ;
        RECT  6.50 4.10 7.00 8.10 ;
        RECT  7.00 7.60 7.50 10.55 ;
        RECT  7.00 8.90 7.70 10.55 ;
        RECT  6.50 4.10 8.15 5.00 ;
        RECT  4.50 7.60 10.20 8.10 ;
        RECT  9.70 7.60 10.20 10.55 ;
        RECT  9.70 8.95 10.40 10.55 ;
        RECT  13.75 2.45 14.25 4.80 ;
        RECT  6.50 4.10 14.25 4.80 ;
        RECT  13.75 2.45 15.05 3.15 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  21.25 5.25 22.15 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  22.65 5.40 23.55 6.30 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  19.15 4.45 19.65 6.30 ;
        RECT  18.45 5.40 19.65 6.30 ;
        RECT  19.15 4.45 19.85 5.15 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.10 17.95 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.30 2.55 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  0.25 4.10 1.15 5.00 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.80 8.30 3.50 11.00 ;
        RECT  5.65 8.55 6.35 11.00 ;
        RECT  8.35 8.55 9.05 11.00 ;
        RECT  11.05 8.35 11.75 11.00 ;
        RECT  12.55 9.20 14.15 11.00 ;
        RECT  20.05 8.20 20.75 11.00 ;
        RECT  0.00 11.00 23.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.45 2.00 1.15 3.65 ;
        RECT  3.30 2.00 4.00 3.70 ;
        RECT  17.25 2.00 17.95 3.05 ;
        RECT  19.95 2.00 20.65 3.10 ;
        RECT  22.65 2.00 23.35 3.10 ;
        RECT  0.00 0.00 23.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.65 6.75 1.15 10.55 ;
        RECT  0.45 8.50 1.15 10.55 ;
        RECT  1.80 2.95 2.50 3.65 ;
        RECT  2.00 2.95 2.50 4.85 ;
        RECT  2.00 4.35 3.50 4.85 ;
        RECT  3.00 4.35 3.50 7.25 ;
        RECT  0.65 6.75 3.50 7.25 ;
        RECT  3.00 6.25 4.45 6.95 ;
        RECT  0.65 6.75 4.45 6.95 ;
        RECT  7.65 5.50 8.15 7.15 ;
        RECT  7.45 6.45 8.15 7.15 ;
        RECT  10.15 6.45 10.85 7.15 ;
        RECT  10.15 6.65 13.75 7.15 ;
        RECT  13.25 6.65 13.75 8.65 ;
        RECT  7.65 5.50 15.20 6.00 ;
        RECT  13.25 8.15 15.35 8.65 ;
        RECT  14.70 3.60 15.20 7.60 ;
        RECT  14.85 8.15 15.35 10.55 ;
        RECT  15.90 2.45 16.60 4.10 ;
        RECT  14.70 3.60 16.60 4.10 ;
        RECT  14.70 7.10 17.40 7.60 ;
        RECT  16.70 7.10 17.40 9.15 ;
        RECT  15.80 8.45 17.40 9.15 ;
        RECT  15.90 3.50 19.10 4.00 ;
        RECT  18.60 2.45 19.10 4.00 ;
        RECT  14.70 3.60 19.10 4.00 ;
        RECT  18.60 2.45 19.30 3.15 ;
        RECT  19.00 7.15 19.50 10.55 ;
        RECT  14.85 10.05 19.50 10.55 ;
        RECT  20.30 4.30 20.80 7.65 ;
        RECT  21.30 2.45 21.80 4.80 ;
        RECT  20.30 4.30 21.80 4.80 ;
        RECT  21.30 2.45 22.00 3.15 ;
        RECT  19.00 7.15 23.25 7.65 ;
        RECT  22.55 7.15 23.25 10.55 ;
    END
END OR7X4
MACRO OR8X1
    CLASS CORE ;
    FOREIGN OR8X1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  7.20 4.50 7.45 10.20 ;
        RECT  6.75 7.70 7.45 10.20 ;
        RECT  7.20 4.50 7.70 8.20 ;
        RECT  6.75 7.70 10.15 8.20 ;
        RECT  8.75 2.45 9.45 5.00 ;
        RECT  8.65 4.10 9.55 5.00 ;
        RECT  7.20 4.50 9.55 5.00 ;
        RECT  9.45 7.70 10.15 10.20 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.25 17.95 6.30 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.40 19.35 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  14.25 4.10 15.15 5.00 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  12.85 4.10 13.75 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  11.45 4.10 12.35 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.40 5.50 6.30 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  5.40 8.65 6.10 11.00 ;
        RECT  8.10 8.65 8.80 11.00 ;
        RECT  15.85 8.20 16.55 11.00 ;
        RECT  0.00 11.00 19.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.55 2.00 3.25 3.65 ;
        RECT  5.40 2.00 6.10 3.65 ;
        RECT  12.90 2.00 13.60 2.70 ;
        RECT  15.75 2.00 16.45 3.10 ;
        RECT  18.45 2.00 19.15 3.15 ;
        RECT  0.00 0.00 19.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.45 8.05 1.15 10.55 ;
        RECT  1.20 2.95 1.90 3.65 ;
        RECT  1.40 2.95 1.90 4.70 ;
        RECT  2.25 6.75 2.75 8.75 ;
        RECT  0.45 8.05 2.75 8.75 ;
        RECT  3.90 2.95 4.40 4.70 ;
        RECT  3.90 2.95 4.60 3.65 ;
        RECT  1.40 4.20 6.45 4.70 ;
        RECT  5.95 4.20 6.45 7.25 ;
        RECT  2.25 6.75 6.45 7.25 ;
        RECT  5.95 4.90 6.75 5.60 ;
        RECT  8.35 6.05 8.85 7.25 ;
        RECT  8.15 6.55 8.85 7.25 ;
        RECT  10.50 3.15 11.00 6.55 ;
        RECT  10.70 7.00 11.15 10.55 ;
        RECT  10.65 7.45 11.15 10.55 ;
        RECT  10.70 7.00 11.40 7.70 ;
        RECT  10.65 7.45 11.40 7.70 ;
        RECT  11.40 2.45 12.10 3.65 ;
        RECT  8.35 6.05 13.00 6.55 ;
        RECT  12.50 6.05 13.00 9.15 ;
        RECT  12.50 7.10 13.20 9.15 ;
        RECT  11.60 8.45 13.20 9.15 ;
        RECT  14.40 2.45 15.10 3.65 ;
        RECT  10.50 3.15 15.10 3.65 ;
        RECT  14.80 7.15 15.30 10.55 ;
        RECT  10.65 10.05 15.30 10.55 ;
        RECT  16.00 4.30 16.50 7.65 ;
        RECT  17.10 2.45 17.60 4.80 ;
        RECT  16.00 4.30 17.60 4.80 ;
        RECT  17.10 2.45 17.80 3.15 ;
        RECT  14.80 7.15 19.05 7.65 ;
        RECT  18.35 7.15 19.05 10.55 ;
    END
END OR8X1
MACRO OR8X2
    CLASS CORE ;
    FOREIGN OR8X2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 22.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  7.80 4.50 8.30 10.20 ;
        RECT  7.75 7.70 8.45 10.20 ;
        RECT  8.65 4.10 9.55 5.00 ;
        RECT  7.60 7.70 11.15 8.20 ;
        RECT  10.45 7.70 11.15 10.20 ;
        RECT  8.65 4.25 12.85 5.00 ;
        RECT  12.15 2.45 12.85 5.00 ;
        RECT  7.80 4.50 12.85 5.00 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.25 20.75 6.30 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  21.25 5.40 22.15 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  17.05 4.10 17.95 5.00 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  15.65 4.10 16.55 5.00 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  14.25 4.10 15.15 5.00 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  5.85 4.10 6.75 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  4.45 5.30 5.35 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  6.25 7.70 6.95 11.00 ;
        RECT  9.10 8.65 9.80 11.00 ;
        RECT  12.00 8.30 12.70 11.00 ;
        RECT  18.65 8.20 19.35 11.00 ;
        RECT  0.00 11.00 22.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  2.55 2.00 3.25 3.65 ;
        RECT  5.25 2.00 5.95 3.65 ;
        RECT  6.75 2.00 7.45 3.65 ;
        RECT  15.70 2.00 16.40 2.70 ;
        RECT  18.55 2.00 19.25 3.10 ;
        RECT  21.25 2.00 21.95 3.15 ;
        RECT  0.00 0.00 22.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.20 2.95 1.90 3.65 ;
        RECT  1.40 2.95 1.90 4.70 ;
        RECT  1.30 8.05 2.00 10.55 ;
        RECT  3.10 6.75 3.60 8.75 ;
        RECT  3.50 4.20 3.60 8.75 ;
        RECT  1.30 8.05 3.60 8.75 ;
        RECT  3.90 2.95 4.00 7.25 ;
        RECT  3.50 4.20 4.00 7.25 ;
        RECT  3.90 2.95 4.40 4.70 ;
        RECT  1.40 4.20 4.40 4.70 ;
        RECT  3.90 2.95 4.60 3.65 ;
        RECT  6.65 6.10 7.15 7.25 ;
        RECT  3.10 6.75 7.15 7.25 ;
        RECT  6.65 6.10 7.35 6.80 ;
        RECT  3.10 6.75 7.35 6.80 ;
        RECT  8.95 6.05 9.45 7.25 ;
        RECT  8.75 6.55 9.45 7.25 ;
        RECT  11.60 7.00 12.30 7.70 ;
        RECT  11.60 7.20 13.90 7.70 ;
        RECT  13.30 3.15 13.80 6.55 ;
        RECT  13.40 7.20 13.90 10.55 ;
        RECT  14.20 2.45 14.90 3.65 ;
        RECT  8.95 6.05 15.80 6.55 ;
        RECT  15.30 6.05 15.80 9.15 ;
        RECT  15.30 7.10 16.00 9.15 ;
        RECT  14.40 8.45 16.00 9.15 ;
        RECT  17.20 2.45 17.90 3.65 ;
        RECT  13.30 3.15 17.90 3.65 ;
        RECT  17.60 7.15 18.10 10.55 ;
        RECT  13.40 10.05 18.10 10.55 ;
        RECT  18.80 4.30 19.30 7.65 ;
        RECT  19.90 2.45 20.40 4.80 ;
        RECT  18.80 4.30 20.40 4.80 ;
        RECT  19.90 2.45 20.60 3.15 ;
        RECT  17.60 7.15 21.85 7.65 ;
        RECT  21.15 7.15 21.85 10.55 ;
    END
END OR8X2
MACRO OR8X3
    CLASS CORE ;
    FOREIGN OR8X3 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 23.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  7.10 7.40 7.80 10.55 ;
        RECT  9.85 4.10 10.35 10.55 ;
        RECT  9.80 7.40 10.50 10.55 ;
        RECT  9.85 4.10 10.95 5.00 ;
        RECT  7.10 7.40 13.20 7.90 ;
        RECT  12.50 7.40 13.20 10.55 ;
        RECT  13.75 2.45 14.25 4.80 ;
        RECT  9.45 4.10 14.25 4.80 ;
        RECT  13.75 2.45 15.05 3.15 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  21.25 5.25 22.15 6.30 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  22.65 5.40 23.55 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  19.15 4.45 19.65 6.30 ;
        RECT  18.45 5.40 19.65 6.30 ;
        RECT  19.15 4.45 19.85 5.15 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  17.05 5.10 17.95 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  15.65 5.40 16.55 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  4.45 4.10 5.35 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.30 3.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  5.55 7.70 6.25 11.00 ;
        RECT  8.45 8.35 9.15 11.00 ;
        RECT  11.15 8.35 11.85 11.00 ;
        RECT  13.85 8.35 14.55 11.00 ;
        RECT  20.05 8.20 20.75 11.00 ;
        RECT  0.00 11.00 23.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.90 2.00 2.60 3.65 ;
        RECT  4.60 2.00 5.30 3.65 ;
        RECT  6.10 2.00 6.80 3.65 ;
        RECT  17.25 2.00 17.95 3.05 ;
        RECT  19.95 2.00 20.65 3.10 ;
        RECT  22.65 2.00 23.35 3.10 ;
        RECT  0.00 0.00 23.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.55 2.95 1.25 3.65 ;
        RECT  0.50 8.05 1.20 10.55 ;
        RECT  0.75 2.95 1.25 4.70 ;
        RECT  2.10 4.20 2.60 8.75 ;
        RECT  0.50 8.05 2.90 8.75 ;
        RECT  3.25 2.95 3.75 4.70 ;
        RECT  0.75 4.20 3.75 4.70 ;
        RECT  3.25 2.95 3.95 3.65 ;
        RECT  6.15 6.25 6.65 7.25 ;
        RECT  2.10 6.75 6.65 7.25 ;
        RECT  6.15 6.25 7.25 6.95 ;
        RECT  2.10 6.75 7.25 6.95 ;
        RECT  10.80 6.25 11.50 6.95 ;
        RECT  14.70 3.60 15.20 7.25 ;
        RECT  10.80 6.25 15.20 6.75 ;
        RECT  15.00 9.85 15.70 10.55 ;
        RECT  15.90 2.45 16.60 4.10 ;
        RECT  14.70 3.60 16.60 4.10 ;
        RECT  14.70 6.75 17.40 7.25 ;
        RECT  16.70 6.75 17.40 9.15 ;
        RECT  15.80 8.45 17.40 9.15 ;
        RECT  15.90 3.50 19.10 4.00 ;
        RECT  18.60 2.45 19.10 4.00 ;
        RECT  14.70 3.60 19.10 4.00 ;
        RECT  18.60 2.45 19.30 3.15 ;
        RECT  19.00 7.15 19.50 10.55 ;
        RECT  15.00 10.05 19.50 10.55 ;
        RECT  20.30 4.30 20.80 7.65 ;
        RECT  21.30 2.45 21.80 4.80 ;
        RECT  20.30 4.30 21.80 4.80 ;
        RECT  21.30 2.45 22.00 3.15 ;
        RECT  19.00 7.15 23.25 7.65 ;
        RECT  22.55 7.15 23.25 10.55 ;
    END
END OR8X3
MACRO OR8X4
    CLASS CORE ;
    FOREIGN OR8X4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 26.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  7.30 7.60 7.80 10.55 ;
        RECT  7.10 8.90 7.80 10.55 ;
        RECT  9.30 4.10 9.80 8.10 ;
        RECT  9.80 7.60 10.30 10.55 ;
        RECT  9.80 8.90 10.50 10.55 ;
        RECT  9.30 4.10 10.95 5.00 ;
        RECT  7.30 7.60 13.00 8.10 ;
        RECT  12.50 7.60 13.00 10.55 ;
        RECT  12.50 8.95 13.20 10.55 ;
        RECT  16.55 2.45 17.05 4.80 ;
        RECT  9.30 4.10 17.05 4.80 ;
        RECT  16.55 2.45 17.85 3.15 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  24.05 5.25 24.95 6.30 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.75 ;
        PORT
        LAYER M1M ;
        RECT  25.45 5.40 26.35 6.30 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  21.95 4.45 22.45 6.30 ;
        RECT  21.25 5.40 22.45 6.30 ;
        RECT  21.95 4.45 22.65 5.15 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  19.85 5.10 20.75 6.30 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  18.45 5.40 19.35 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  4.45 4.10 5.35 5.00 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.30 3.95 6.30 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  0.25 5.40 1.15 6.30 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  5.70 8.15 6.40 11.00 ;
        RECT  8.45 8.55 9.15 11.00 ;
        RECT  11.15 8.55 11.85 11.00 ;
        RECT  13.85 8.35 14.55 11.00 ;
        RECT  15.35 9.20 16.95 11.00 ;
        RECT  22.85 8.20 23.55 11.00 ;
        RECT  0.00 11.00 26.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.90 2.00 2.60 3.65 ;
        RECT  4.60 2.00 5.30 3.65 ;
        RECT  6.10 2.00 6.80 5.30 ;
        RECT  20.05 2.00 20.75 3.05 ;
        RECT  22.75 2.00 23.45 3.10 ;
        RECT  25.45 2.00 26.15 3.10 ;
        RECT  0.00 0.00 26.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.55 2.95 1.25 3.65 ;
        RECT  0.45 8.05 1.15 10.55 ;
        RECT  0.75 2.95 1.25 4.70 ;
        RECT  2.05 4.20 2.55 8.75 ;
        RECT  0.45 8.05 2.95 8.75 ;
        RECT  3.25 2.95 3.75 4.70 ;
        RECT  0.75 4.20 3.75 4.70 ;
        RECT  3.25 2.95 3.95 3.65 ;
        RECT  6.50 6.25 7.00 7.25 ;
        RECT  2.05 6.75 7.00 7.25 ;
        RECT  6.50 6.25 7.25 6.95 ;
        RECT  2.05 6.75 7.25 6.95 ;
        RECT  10.45 5.50 10.95 7.15 ;
        RECT  10.25 6.45 10.95 7.15 ;
        RECT  12.95 6.45 13.65 7.15 ;
        RECT  12.95 6.65 16.55 7.15 ;
        RECT  16.05 6.65 16.55 8.65 ;
        RECT  10.45 5.50 18.00 6.00 ;
        RECT  16.05 8.15 18.15 8.65 ;
        RECT  17.50 3.60 18.00 7.60 ;
        RECT  17.65 8.15 18.15 10.55 ;
        RECT  18.70 2.45 19.40 4.10 ;
        RECT  17.50 3.60 19.40 4.10 ;
        RECT  17.50 7.10 20.20 7.60 ;
        RECT  19.50 7.10 20.20 9.15 ;
        RECT  18.60 8.45 20.20 9.15 ;
        RECT  18.70 3.50 21.90 4.00 ;
        RECT  21.40 2.45 21.90 4.00 ;
        RECT  17.50 3.60 21.90 4.00 ;
        RECT  21.40 2.45 22.10 3.15 ;
        RECT  21.80 7.15 22.30 10.55 ;
        RECT  17.65 10.05 22.30 10.55 ;
        RECT  23.10 4.30 23.60 7.65 ;
        RECT  24.10 2.45 24.60 4.80 ;
        RECT  23.10 4.30 24.60 4.80 ;
        RECT  24.10 2.45 24.80 3.15 ;
        RECT  21.80 7.15 26.05 7.65 ;
        RECT  25.35 7.15 26.05 10.55 ;
    END
END OR8X4
MACRO SDFFRSX1
    CLASS CORE ;
    FOREIGN SDFFRSX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 35.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  16.80 2.55 17.95 3.45 ;
        RECT  17.05 2.55 17.95 3.75 ;
        RECT  16.80 2.55 29.50 3.05 ;
        RECT  28.80 2.55 29.50 3.25 ;
        END
    END SN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  1.45 5.60 2.55 6.30 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END SD
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  20.45 5.75 21.15 6.45 ;
        RECT  22.65 5.35 23.55 6.35 ;
        RECT  20.45 5.85 23.55 6.35 ;
        RECT  22.65 5.50 24.90 6.20 ;
        RECT  20.45 5.85 24.90 6.20 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  31.15 2.65 31.85 4.30 ;
        RECT  31.15 7.25 31.85 9.75 ;
        RECT  31.15 3.80 32.95 4.30 ;
        RECT  32.45 3.80 32.95 7.75 ;
        RECT  31.15 7.25 32.95 7.75 ;
        RECT  32.45 5.35 33.35 6.35 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  33.85 2.65 34.55 3.35 ;
        RECT  34.05 2.65 34.55 9.75 ;
        RECT  33.85 7.95 34.55 9.75 ;
        RECT  33.75 7.95 34.75 8.95 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  6.50 8.10 7.20 11.00 ;
        RECT  10.75 8.85 11.45 11.00 ;
        RECT  16.80 8.45 17.50 11.00 ;
        RECT  19.65 7.30 20.35 11.00 ;
        RECT  19.65 7.30 25.35 7.80 ;
        RECT  24.65 7.30 25.35 8.35 ;
        RECT  26.85 9.25 27.55 11.00 ;
        RECT  29.55 9.25 30.25 11.00 ;
        RECT  32.50 8.25 33.20 11.00 ;
        RECT  0.00 11.00 35.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.45 ;
        RECT  6.50 2.00 7.20 4.40 ;
        RECT  10.70 2.00 11.40 3.95 ;
        RECT  15.85 2.00 16.35 5.00 ;
        RECT  17.00 4.50 17.70 5.20 ;
        RECT  18.55 3.55 19.05 5.00 ;
        RECT  15.85 4.50 19.05 5.00 ;
        RECT  18.55 3.55 21.85 4.05 ;
        RECT  21.15 3.55 21.85 4.25 ;
        RECT  26.85 3.55 27.55 4.25 ;
        RECT  26.85 3.75 30.65 4.25 ;
        RECT  30.15 2.00 30.65 5.50 ;
        RECT  30.15 4.80 31.40 5.50 ;
        RECT  32.50 2.00 33.20 3.30 ;
        RECT  0.00 0.00 35.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.15 3.95 5.20 4.45 ;
        RECT  0.45 3.75 0.95 9.90 ;
        RECT  0.45 3.75 1.15 4.45 ;
        RECT  0.45 8.10 1.15 9.90 ;
        RECT  3.50 6.85 4.20 7.55 ;
        RECT  0.45 7.05 4.20 7.55 ;
        RECT  4.70 3.75 4.85 9.90 ;
        RECT  4.15 8.15 4.85 9.90 ;
        RECT  4.70 3.75 5.05 8.65 ;
        RECT  4.15 3.75 5.05 4.45 ;
        RECT  4.70 3.95 5.20 8.65 ;
        RECT  4.15 8.15 5.20 8.65 ;
        RECT  7.85 3.80 8.55 4.95 ;
        RECT  7.85 7.70 8.55 9.85 ;
        RECT  7.85 4.45 9.30 4.95 ;
        RECT  7.85 7.70 9.25 8.40 ;
        RECT  8.60 4.45 9.30 5.55 ;
        RECT  9.35 3.25 10.25 3.95 ;
        RECT  9.45 6.40 10.15 7.25 ;
        RECT  4.70 6.75 10.15 7.25 ;
        RECT  9.75 3.25 10.25 5.20 ;
        RECT  9.80 7.90 10.30 9.85 ;
        RECT  9.35 9.15 10.30 9.85 ;
        RECT  9.75 4.70 11.10 5.20 ;
        RECT  10.60 4.70 11.10 8.40 ;
        RECT  9.80 7.90 11.10 8.40 ;
        RECT  10.60 6.05 13.15 6.55 ;
        RECT  12.45 6.05 13.15 6.75 ;
        RECT  13.45 4.80 14.15 5.50 ;
        RECT  13.65 4.80 14.15 7.55 ;
        RECT  13.65 6.85 14.40 7.55 ;
        RECT  13.10 3.20 15.35 3.90 ;
        RECT  14.85 3.20 15.35 9.40 ;
        RECT  13.25 8.70 15.35 9.40 ;
        RECT  16.35 5.65 17.05 6.35 ;
        RECT  17.50 6.90 18.20 7.60 ;
        RECT  14.85 7.10 18.20 7.60 ;
        RECT  18.65 5.65 19.15 9.15 ;
        RECT  18.15 8.45 19.15 9.15 ;
        RECT  19.50 4.55 20.00 6.15 ;
        RECT  16.35 5.65 20.00 6.15 ;
        RECT  19.50 4.55 20.20 5.25 ;
        RECT  22.00 8.30 22.70 10.05 ;
        RECT  23.50 3.55 24.20 4.25 ;
        RECT  24.50 8.85 25.20 9.95 ;
        RECT  23.50 3.75 26.35 4.25 ;
        RECT  25.85 3.75 26.35 9.35 ;
        RECT  22.00 8.85 26.35 9.35 ;
        RECT  26.85 4.75 29.05 5.45 ;
        RECT  28.20 8.25 28.90 9.90 ;
        RECT  28.55 4.75 29.05 6.55 ;
        RECT  28.95 7.05 29.65 7.75 ;
        RECT  25.85 7.25 29.65 7.75 ;
        RECT  30.15 6.05 30.65 8.75 ;
        RECT  28.20 8.25 30.65 8.75 ;
        RECT  28.55 6.05 31.95 6.55 ;
        RECT  31.25 6.05 31.95 6.75 ;
    END
END SDFFRSX1
MACRO SDFFRSX2
    CLASS CORE ;
    FOREIGN SDFFRSX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 35.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  16.80 2.55 17.95 3.45 ;
        RECT  17.05 2.55 17.95 3.75 ;
        RECT  16.80 2.55 29.50 3.05 ;
        RECT  28.80 2.55 29.50 3.25 ;
        END
    END SN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  1.45 5.60 2.55 6.30 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END SD
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  20.45 5.75 21.15 6.45 ;
        RECT  22.65 5.35 23.55 6.35 ;
        RECT  20.45 5.85 23.55 6.35 ;
        RECT  22.65 5.50 24.90 6.20 ;
        RECT  20.45 5.85 24.90 6.20 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  33.85 2.65 34.55 3.35 ;
        RECT  34.05 2.65 34.55 10.50 ;
        RECT  33.85 7.95 34.55 10.50 ;
        RECT  33.75 7.95 34.75 8.95 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END CN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  31.15 2.65 31.85 4.30 ;
        RECT  31.15 7.25 31.85 10.50 ;
        RECT  31.15 3.80 32.95 4.30 ;
        RECT  32.45 3.80 32.95 7.75 ;
        RECT  31.15 7.25 32.95 7.75 ;
        RECT  32.45 5.35 33.35 6.35 ;
        END
    END QN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  6.50 8.10 7.20 11.00 ;
        RECT  10.75 8.85 11.45 11.00 ;
        RECT  16.80 8.45 17.50 11.00 ;
        RECT  19.65 7.30 20.35 11.00 ;
        RECT  19.65 7.30 25.35 7.80 ;
        RECT  24.65 7.30 25.35 8.35 ;
        RECT  26.85 9.25 27.55 11.00 ;
        RECT  29.55 9.25 30.25 11.00 ;
        RECT  32.50 8.25 33.20 11.00 ;
        RECT  0.00 11.00 35.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.45 ;
        RECT  6.50 2.00 7.20 4.40 ;
        RECT  10.70 2.00 11.40 3.95 ;
        RECT  15.85 2.00 16.35 5.00 ;
        RECT  17.00 4.50 17.70 5.20 ;
        RECT  18.55 3.55 19.05 5.00 ;
        RECT  15.85 4.50 19.05 5.00 ;
        RECT  18.55 3.55 21.85 4.05 ;
        RECT  21.15 3.55 21.85 4.25 ;
        RECT  26.85 3.55 27.55 4.25 ;
        RECT  26.85 3.75 30.65 4.25 ;
        RECT  30.15 2.00 30.65 5.50 ;
        RECT  30.15 4.80 31.40 5.50 ;
        RECT  32.50 2.00 33.20 3.30 ;
        RECT  0.00 0.00 35.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.15 3.95 5.20 4.45 ;
        RECT  0.45 3.75 0.95 9.90 ;
        RECT  0.45 3.75 1.15 4.45 ;
        RECT  0.45 8.10 1.15 9.90 ;
        RECT  3.50 6.85 4.20 7.55 ;
        RECT  0.45 7.05 4.20 7.55 ;
        RECT  4.70 3.75 4.85 9.90 ;
        RECT  4.15 8.15 4.85 9.90 ;
        RECT  4.70 3.75 5.05 8.65 ;
        RECT  4.15 3.75 5.05 4.45 ;
        RECT  4.70 3.95 5.20 8.65 ;
        RECT  4.15 8.15 5.20 8.65 ;
        RECT  7.85 3.80 8.55 4.95 ;
        RECT  7.85 7.70 8.55 9.85 ;
        RECT  7.85 4.45 9.30 4.95 ;
        RECT  7.85 7.70 9.25 8.40 ;
        RECT  8.60 4.45 9.30 5.55 ;
        RECT  9.35 3.25 10.25 3.95 ;
        RECT  9.45 6.40 10.15 7.25 ;
        RECT  4.70 6.75 10.15 7.25 ;
        RECT  9.75 3.25 10.25 5.20 ;
        RECT  9.80 7.90 10.30 9.85 ;
        RECT  9.35 9.15 10.30 9.85 ;
        RECT  9.75 4.70 11.10 5.20 ;
        RECT  10.60 4.70 11.10 8.40 ;
        RECT  9.80 7.90 11.10 8.40 ;
        RECT  10.60 6.05 13.15 6.55 ;
        RECT  12.45 6.05 13.15 6.75 ;
        RECT  13.45 4.80 14.15 5.50 ;
        RECT  13.65 4.80 14.15 7.55 ;
        RECT  13.65 6.85 14.40 7.55 ;
        RECT  13.10 3.20 15.35 3.90 ;
        RECT  14.85 3.20 15.35 9.40 ;
        RECT  13.25 8.70 15.35 9.40 ;
        RECT  16.35 5.65 17.05 6.35 ;
        RECT  17.50 6.90 18.20 7.60 ;
        RECT  14.85 7.10 18.20 7.60 ;
        RECT  18.65 5.65 19.15 9.15 ;
        RECT  18.15 8.45 19.15 9.15 ;
        RECT  19.50 4.55 20.00 6.15 ;
        RECT  16.35 5.65 20.00 6.15 ;
        RECT  19.50 4.55 20.20 5.25 ;
        RECT  22.00 8.30 22.70 10.05 ;
        RECT  23.50 3.55 24.20 4.25 ;
        RECT  24.50 8.85 25.20 9.95 ;
        RECT  23.50 3.75 26.35 4.25 ;
        RECT  25.85 3.75 26.35 9.35 ;
        RECT  22.00 8.85 26.35 9.35 ;
        RECT  26.85 4.75 29.05 5.45 ;
        RECT  28.20 8.25 28.90 9.90 ;
        RECT  28.55 4.75 29.05 6.55 ;
        RECT  28.95 7.05 29.65 7.75 ;
        RECT  25.85 7.25 29.65 7.75 ;
        RECT  30.15 6.05 30.65 8.75 ;
        RECT  28.20 8.25 30.65 8.75 ;
        RECT  28.55 6.05 31.95 6.55 ;
        RECT  31.25 6.05 31.95 6.75 ;
    END
END SDFFRSX2
MACRO SDFFRSX4
    CLASS CORE ;
    FOREIGN SDFFRSX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 37.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  16.80 2.55 17.95 3.45 ;
        RECT  17.05 2.55 17.95 3.75 ;
        RECT  16.80 2.55 29.50 3.05 ;
        RECT  28.80 2.55 29.50 3.25 ;
        END
    END SN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  1.45 5.60 2.55 6.30 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END SD
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  20.45 5.75 21.15 6.45 ;
        RECT  22.65 5.35 23.55 6.35 ;
        RECT  20.45 5.85 23.55 6.35 ;
        RECT  22.65 5.50 24.90 6.20 ;
        RECT  20.45 5.85 24.90 6.20 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  35.30 2.50 36.00 4.10 ;
        RECT  35.50 2.50 36.00 10.50 ;
        RECT  35.30 5.35 36.00 10.50 ;
        RECT  35.15 5.35 36.15 6.35 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END CN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  32.60 2.50 33.10 10.50 ;
        RECT  32.60 2.50 33.30 4.10 ;
        RECT  32.60 8.10 33.30 10.50 ;
        RECT  32.45 5.35 33.35 6.35 ;
        END
    END QN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  6.50 8.10 7.20 11.00 ;
        RECT  10.75 8.85 11.45 11.00 ;
        RECT  16.80 8.45 17.50 11.00 ;
        RECT  19.65 7.30 20.35 11.00 ;
        RECT  19.65 7.30 25.35 7.80 ;
        RECT  24.65 7.30 25.35 8.35 ;
        RECT  26.85 9.25 27.55 11.00 ;
        RECT  29.55 9.25 30.25 11.00 ;
        RECT  31.25 8.10 31.95 11.00 ;
        RECT  33.95 8.10 34.65 11.00 ;
        RECT  36.65 8.10 37.35 11.00 ;
        RECT  0.00 11.00 37.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.45 ;
        RECT  6.50 2.00 7.20 4.40 ;
        RECT  10.70 2.00 11.40 3.95 ;
        RECT  15.85 2.00 16.35 5.00 ;
        RECT  17.00 4.50 17.70 5.20 ;
        RECT  18.55 3.55 19.05 5.00 ;
        RECT  15.85 4.50 19.05 5.00 ;
        RECT  18.55 3.55 21.85 4.05 ;
        RECT  21.15 3.55 21.85 4.25 ;
        RECT  26.85 3.55 27.55 4.25 ;
        RECT  26.85 3.75 30.65 4.25 ;
        RECT  30.15 2.00 30.65 5.50 ;
        RECT  30.15 4.80 31.40 5.50 ;
        RECT  31.10 2.00 31.80 3.90 ;
        RECT  33.95 2.00 34.65 4.10 ;
        RECT  36.65 2.00 37.35 4.10 ;
        RECT  0.00 0.00 37.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.15 3.95 5.20 4.45 ;
        RECT  0.45 3.75 0.95 9.90 ;
        RECT  0.45 3.75 1.15 4.45 ;
        RECT  0.45 8.10 1.15 9.90 ;
        RECT  3.50 6.85 4.20 7.55 ;
        RECT  0.45 7.05 4.20 7.55 ;
        RECT  4.70 3.75 4.85 9.90 ;
        RECT  4.15 8.15 4.85 9.90 ;
        RECT  4.70 3.75 5.05 8.65 ;
        RECT  4.15 3.75 5.05 4.45 ;
        RECT  4.70 3.95 5.20 8.65 ;
        RECT  4.15 8.15 5.20 8.65 ;
        RECT  7.85 3.80 8.55 4.95 ;
        RECT  7.85 7.70 8.55 9.85 ;
        RECT  7.85 4.45 9.30 4.95 ;
        RECT  7.85 7.70 9.25 8.40 ;
        RECT  8.60 4.45 9.30 5.55 ;
        RECT  9.35 3.25 10.25 3.95 ;
        RECT  9.45 6.40 10.15 7.25 ;
        RECT  4.70 6.75 10.15 7.25 ;
        RECT  9.75 3.25 10.25 5.20 ;
        RECT  9.80 7.90 10.30 9.85 ;
        RECT  9.35 9.15 10.30 9.85 ;
        RECT  9.75 4.70 11.10 5.20 ;
        RECT  10.60 4.70 11.10 8.40 ;
        RECT  9.80 7.90 11.10 8.40 ;
        RECT  10.60 6.05 13.15 6.55 ;
        RECT  12.45 6.05 13.15 6.75 ;
        RECT  13.45 4.80 14.15 5.50 ;
        RECT  13.65 4.80 14.15 7.55 ;
        RECT  13.65 6.85 14.40 7.55 ;
        RECT  13.10 3.20 15.35 3.90 ;
        RECT  14.85 3.20 15.35 9.40 ;
        RECT  13.25 8.70 15.35 9.40 ;
        RECT  16.35 5.65 17.05 6.35 ;
        RECT  17.50 6.90 18.20 7.60 ;
        RECT  14.85 7.10 18.20 7.60 ;
        RECT  18.65 5.65 19.15 9.15 ;
        RECT  18.15 8.45 19.15 9.15 ;
        RECT  19.50 4.55 20.00 6.15 ;
        RECT  16.35 5.65 20.00 6.15 ;
        RECT  19.50 4.55 20.20 5.25 ;
        RECT  22.00 8.30 22.70 10.05 ;
        RECT  23.50 3.55 24.20 4.25 ;
        RECT  24.50 8.85 25.20 9.95 ;
        RECT  23.50 3.75 26.35 4.25 ;
        RECT  25.85 3.75 26.35 9.35 ;
        RECT  22.00 8.85 26.35 9.35 ;
        RECT  26.85 4.75 29.05 5.45 ;
        RECT  28.20 8.25 28.90 9.90 ;
        RECT  28.55 4.75 29.05 6.55 ;
        RECT  28.95 7.05 29.65 7.75 ;
        RECT  25.85 7.25 29.65 7.75 ;
        RECT  30.15 6.05 30.65 8.75 ;
        RECT  28.20 8.25 30.65 8.75 ;
        RECT  28.55 6.05 31.95 6.55 ;
        RECT  31.25 6.05 31.95 6.75 ;
    END
END SDFFRSX4
MACRO SDFFRX1
    CLASS CORE ;
    FOREIGN SDFFRX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 30.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  1.45 5.60 2.55 6.30 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END SD
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  18.45 7.05 19.15 8.40 ;
        RECT  19.85 6.70 20.75 7.60 ;
        RECT  20.25 5.45 20.75 7.60 ;
        RECT  18.45 7.05 20.75 7.60 ;
        RECT  20.90 5.25 21.60 5.95 ;
        RECT  20.25 5.45 21.60 5.95 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  29.65 3.75 30.35 4.45 ;
        RECT  29.85 3.75 30.35 8.85 ;
        RECT  29.65 7.15 30.35 8.85 ;
        RECT  29.65 5.40 30.55 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  26.95 3.75 27.65 4.45 ;
        RECT  27.10 3.75 27.65 8.85 ;
        RECT  26.95 7.15 27.65 8.85 ;
        RECT  26.85 5.40 27.75 6.30 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  6.50 8.10 7.20 11.00 ;
        RECT  10.75 8.85 11.45 11.00 ;
        RECT  15.75 8.35 16.45 11.00 ;
        RECT  19.05 8.90 19.75 11.00 ;
        RECT  24.05 7.40 24.75 11.00 ;
        RECT  28.30 7.15 29.00 11.00 ;
        RECT  24.05 10.70 30.35 11.00 ;
        RECT  0.00 11.00 30.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.45 ;
        RECT  6.50 2.00 7.20 4.40 ;
        RECT  10.70 2.00 11.40 3.95 ;
        RECT  14.75 2.00 16.70 2.40 ;
        RECT  16.00 2.00 16.70 4.60 ;
        RECT  18.20 2.00 18.90 3.25 ;
        RECT  24.05 2.00 24.75 3.95 ;
        RECT  28.30 2.00 29.00 4.45 ;
        RECT  0.00 0.00 30.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.15 3.95 5.20 4.45 ;
        RECT  0.45 3.75 0.95 9.90 ;
        RECT  0.45 3.75 1.15 4.45 ;
        RECT  0.45 8.10 1.15 9.90 ;
        RECT  3.50 6.85 4.20 7.55 ;
        RECT  0.45 7.05 4.20 7.55 ;
        RECT  4.70 3.75 4.85 9.90 ;
        RECT  4.15 8.15 4.85 9.90 ;
        RECT  4.70 3.75 5.05 8.65 ;
        RECT  4.15 3.75 5.05 4.45 ;
        RECT  4.70 3.95 5.20 8.65 ;
        RECT  4.15 8.15 5.20 8.65 ;
        RECT  7.85 3.80 8.55 4.95 ;
        RECT  7.85 7.70 8.55 9.85 ;
        RECT  7.85 4.45 9.30 4.95 ;
        RECT  7.85 7.70 9.25 8.40 ;
        RECT  8.60 4.45 9.30 5.55 ;
        RECT  9.35 3.25 10.25 3.95 ;
        RECT  9.45 6.40 10.15 7.25 ;
        RECT  4.70 6.75 10.15 7.25 ;
        RECT  9.75 3.25 10.25 5.20 ;
        RECT  9.80 7.90 10.30 9.85 ;
        RECT  9.35 9.15 10.30 9.85 ;
        RECT  9.75 4.70 11.10 5.20 ;
        RECT  10.60 4.70 11.10 8.40 ;
        RECT  9.80 7.90 11.10 8.40 ;
        RECT  10.60 6.05 13.15 6.55 ;
        RECT  12.45 6.05 13.15 6.75 ;
        RECT  12.65 7.30 13.35 8.00 ;
        RECT  13.45 4.80 14.15 5.50 ;
        RECT  13.25 8.45 13.95 10.15 ;
        RECT  13.65 4.80 14.15 7.80 ;
        RECT  12.65 7.30 14.15 7.80 ;
        RECT  13.25 3.55 15.10 4.25 ;
        RECT  14.60 3.55 15.10 8.95 ;
        RECT  13.25 8.45 15.10 8.95 ;
        RECT  14.60 6.70 16.95 7.20 ;
        RECT  15.55 5.45 16.25 6.15 ;
        RECT  16.25 6.70 16.95 7.40 ;
        RECT  15.55 5.45 17.95 5.95 ;
        RECT  17.45 4.35 17.95 9.55 ;
        RECT  17.45 8.85 18.25 9.55 ;
        RECT  18.55 4.15 19.25 4.85 ;
        RECT  17.45 4.35 19.25 4.85 ;
        RECT  20.70 3.30 21.40 4.00 ;
        RECT  20.70 3.45 22.60 4.00 ;
        RECT  21.55 7.20 22.10 10.50 ;
        RECT  21.40 8.75 22.10 10.50 ;
        RECT  22.10 3.45 22.60 7.90 ;
        RECT  21.55 7.20 22.60 7.90 ;
        RECT  23.60 4.45 24.30 5.15 ;
        RECT  24.40 5.70 25.10 6.40 ;
        RECT  22.10 5.90 25.10 6.40 ;
        RECT  25.40 3.25 26.10 3.95 ;
        RECT  23.60 4.45 26.10 4.95 ;
        RECT  25.60 3.25 26.10 10.10 ;
        RECT  25.40 7.40 26.10 10.10 ;
    END
END SDFFRX1
MACRO SDFFRX2
    CLASS CORE ;
    FOREIGN SDFFRX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 30.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  1.45 5.60 2.55 6.30 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END SD
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  18.45 7.05 19.15 8.40 ;
        RECT  19.85 6.70 20.75 7.60 ;
        RECT  20.25 5.45 20.75 7.60 ;
        RECT  18.45 7.05 20.75 7.60 ;
        RECT  20.90 5.25 21.60 5.95 ;
        RECT  20.25 5.45 21.60 5.95 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  29.65 2.70 30.35 4.50 ;
        RECT  29.85 2.70 30.35 10.50 ;
        RECT  29.65 7.10 30.35 10.50 ;
        RECT  29.65 5.40 30.55 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  26.95 2.70 27.65 4.50 ;
        RECT  27.10 2.70 27.65 10.50 ;
        RECT  26.95 7.10 27.65 10.50 ;
        RECT  26.85 5.40 27.75 6.30 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  6.50 8.10 7.20 11.00 ;
        RECT  10.75 8.85 11.45 11.00 ;
        RECT  15.75 8.35 16.45 11.00 ;
        RECT  19.05 8.90 19.75 11.00 ;
        RECT  24.05 7.40 24.75 11.00 ;
        RECT  28.30 7.10 29.00 11.00 ;
        RECT  0.00 11.00 30.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.45 ;
        RECT  6.50 2.00 7.20 4.40 ;
        RECT  10.70 2.00 11.40 3.95 ;
        RECT  14.75 2.00 16.70 2.40 ;
        RECT  16.00 2.00 16.70 4.60 ;
        RECT  18.20 2.00 18.90 3.25 ;
        RECT  24.05 2.00 24.75 3.95 ;
        RECT  28.30 2.00 29.00 4.45 ;
        RECT  0.00 0.00 30.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.15 3.95 5.20 4.45 ;
        RECT  0.45 3.75 0.95 9.90 ;
        RECT  0.45 3.75 1.15 4.45 ;
        RECT  0.45 8.10 1.15 9.90 ;
        RECT  3.50 6.85 4.20 7.55 ;
        RECT  0.45 7.05 4.20 7.55 ;
        RECT  4.70 3.75 4.85 9.90 ;
        RECT  4.15 8.15 4.85 9.90 ;
        RECT  4.70 3.75 5.05 8.65 ;
        RECT  4.15 3.75 5.05 4.45 ;
        RECT  4.70 3.95 5.20 8.65 ;
        RECT  4.15 8.15 5.20 8.65 ;
        RECT  7.85 3.80 8.55 4.95 ;
        RECT  7.85 7.70 8.55 9.85 ;
        RECT  7.85 4.45 9.30 4.95 ;
        RECT  7.85 7.70 9.25 8.40 ;
        RECT  8.60 4.45 9.30 5.55 ;
        RECT  9.35 3.25 10.25 3.95 ;
        RECT  9.45 6.40 10.15 7.25 ;
        RECT  4.70 6.75 10.15 7.25 ;
        RECT  9.75 3.25 10.25 5.20 ;
        RECT  9.80 7.90 10.30 9.85 ;
        RECT  9.35 9.15 10.30 9.85 ;
        RECT  9.75 4.70 11.10 5.20 ;
        RECT  10.60 4.70 11.10 8.40 ;
        RECT  9.80 7.90 11.10 8.40 ;
        RECT  10.60 6.05 13.15 6.55 ;
        RECT  12.45 6.05 13.15 6.75 ;
        RECT  12.65 7.30 13.35 8.00 ;
        RECT  13.45 4.80 14.15 5.50 ;
        RECT  13.25 8.45 13.95 10.15 ;
        RECT  13.65 4.80 14.15 7.80 ;
        RECT  12.65 7.30 14.15 7.80 ;
        RECT  13.25 3.55 15.10 4.25 ;
        RECT  14.60 3.55 15.10 8.95 ;
        RECT  13.25 8.45 15.10 8.95 ;
        RECT  14.60 6.70 16.95 7.20 ;
        RECT  15.55 5.45 16.25 6.15 ;
        RECT  16.25 6.70 16.95 7.40 ;
        RECT  15.55 5.45 17.95 5.95 ;
        RECT  17.45 4.35 17.95 9.55 ;
        RECT  17.45 8.85 18.25 9.55 ;
        RECT  18.55 4.15 19.25 4.85 ;
        RECT  17.45 4.35 19.25 4.85 ;
        RECT  20.70 3.30 21.40 4.00 ;
        RECT  20.70 3.45 22.60 4.00 ;
        RECT  21.55 7.20 22.10 10.50 ;
        RECT  21.40 8.75 22.10 10.50 ;
        RECT  22.10 3.45 22.60 7.90 ;
        RECT  21.55 7.20 22.60 7.90 ;
        RECT  23.60 4.45 24.30 5.15 ;
        RECT  24.40 5.70 25.10 6.40 ;
        RECT  22.10 5.90 25.10 6.40 ;
        RECT  25.40 3.25 26.10 3.95 ;
        RECT  23.60 4.45 26.10 4.95 ;
        RECT  25.60 3.25 26.10 10.55 ;
        RECT  25.40 7.40 26.10 10.55 ;
    END
END SDFFRX2
MACRO SDFFRX4
    CLASS CORE ;
    FOREIGN SDFFRX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 33.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  1.45 5.60 2.55 6.30 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END SD
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  18.45 7.05 19.15 8.40 ;
        RECT  19.85 6.70 20.75 7.60 ;
        RECT  20.25 5.45 20.75 7.60 ;
        RECT  18.45 7.05 20.75 7.60 ;
        RECT  20.90 5.25 21.60 5.95 ;
        RECT  20.25 5.45 21.60 5.95 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  31.10 2.50 31.80 4.10 ;
        RECT  31.30 2.50 31.80 10.50 ;
        RECT  31.10 5.35 31.80 10.50 ;
        RECT  30.95 5.35 31.95 6.35 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  28.40 2.50 28.90 10.50 ;
        RECT  28.40 2.50 29.10 4.10 ;
        RECT  28.40 7.10 29.10 10.50 ;
        RECT  28.25 5.35 29.15 6.35 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  6.50 8.10 7.20 11.00 ;
        RECT  10.75 8.85 11.45 11.00 ;
        RECT  15.75 8.35 16.45 11.00 ;
        RECT  19.05 8.90 19.75 11.00 ;
        RECT  24.05 7.40 24.75 11.00 ;
        RECT  27.05 7.10 27.75 11.00 ;
        RECT  29.75 7.10 30.45 11.00 ;
        RECT  32.45 7.10 33.15 11.00 ;
        RECT  0.00 11.00 33.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.45 ;
        RECT  6.50 2.00 7.20 4.40 ;
        RECT  10.70 2.00 11.40 3.95 ;
        RECT  14.75 2.00 16.70 2.40 ;
        RECT  16.00 2.00 16.70 4.60 ;
        RECT  18.20 2.00 18.90 3.25 ;
        RECT  24.05 2.00 24.75 3.95 ;
        RECT  27.05 2.00 27.75 4.10 ;
        RECT  29.75 2.00 30.45 4.10 ;
        RECT  32.45 2.00 33.15 4.10 ;
        RECT  0.00 0.00 33.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.15 3.95 5.20 4.45 ;
        RECT  0.45 3.75 0.95 9.90 ;
        RECT  0.45 3.75 1.15 4.45 ;
        RECT  0.45 8.10 1.15 9.90 ;
        RECT  3.50 6.85 4.20 7.55 ;
        RECT  0.45 7.05 4.20 7.55 ;
        RECT  4.70 3.75 4.85 9.90 ;
        RECT  4.15 8.15 4.85 9.90 ;
        RECT  4.70 3.75 5.05 8.65 ;
        RECT  4.15 3.75 5.05 4.45 ;
        RECT  4.70 3.95 5.20 8.65 ;
        RECT  4.15 8.15 5.20 8.65 ;
        RECT  7.85 3.80 8.55 4.95 ;
        RECT  7.85 7.70 8.55 9.85 ;
        RECT  7.85 4.45 9.30 4.95 ;
        RECT  7.85 7.70 9.25 8.40 ;
        RECT  8.60 4.45 9.30 5.55 ;
        RECT  9.35 3.25 10.25 3.95 ;
        RECT  9.45 6.40 10.15 7.25 ;
        RECT  4.70 6.75 10.15 7.25 ;
        RECT  9.75 3.25 10.25 5.20 ;
        RECT  9.80 7.90 10.30 9.85 ;
        RECT  9.35 9.15 10.30 9.85 ;
        RECT  9.75 4.70 11.10 5.20 ;
        RECT  10.60 4.70 11.10 8.40 ;
        RECT  9.80 7.90 11.10 8.40 ;
        RECT  10.60 6.05 13.15 6.55 ;
        RECT  12.45 6.05 13.15 6.75 ;
        RECT  12.65 7.30 13.35 8.00 ;
        RECT  13.45 4.80 14.15 5.50 ;
        RECT  13.25 8.45 13.95 10.15 ;
        RECT  13.65 4.80 14.15 7.80 ;
        RECT  12.65 7.30 14.15 7.80 ;
        RECT  13.25 3.55 15.10 4.25 ;
        RECT  14.60 3.55 15.10 8.95 ;
        RECT  13.25 8.45 15.10 8.95 ;
        RECT  14.60 6.70 16.95 7.20 ;
        RECT  15.55 5.45 16.25 6.15 ;
        RECT  16.25 6.70 16.95 7.40 ;
        RECT  15.55 5.45 17.95 5.95 ;
        RECT  17.45 4.35 17.95 9.55 ;
        RECT  17.45 8.85 18.25 9.55 ;
        RECT  18.55 4.15 19.25 4.85 ;
        RECT  17.45 4.35 19.25 4.85 ;
        RECT  20.70 3.30 21.40 4.00 ;
        RECT  20.70 3.45 22.60 4.00 ;
        RECT  21.55 7.20 22.10 10.50 ;
        RECT  21.40 8.75 22.10 10.50 ;
        RECT  22.10 3.45 22.60 7.90 ;
        RECT  21.55 7.20 22.60 7.90 ;
        RECT  23.60 4.45 24.30 5.15 ;
        RECT  24.40 5.70 25.10 6.40 ;
        RECT  22.10 5.90 25.10 6.40 ;
        RECT  25.40 3.25 26.10 3.95 ;
        RECT  23.60 4.45 26.10 4.95 ;
        RECT  25.60 3.25 26.10 10.55 ;
        RECT  25.40 7.40 26.10 10.55 ;
    END
END SDFFRX4
MACRO SDFFSX1
    CLASS CORE ;
    FOREIGN SDFFSX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 32.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  16.75 2.55 23.55 3.25 ;
        RECT  22.65 2.55 23.55 3.75 ;
        RECT  16.75 2.55 26.70 3.05 ;
        RECT  26.00 2.55 26.70 3.25 ;
        END
    END SN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  1.45 5.60 2.55 6.30 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END SD
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  28.35 2.65 29.05 4.30 ;
        RECT  28.35 7.25 29.05 9.75 ;
        RECT  28.35 3.80 30.15 4.30 ;
        RECT  29.65 3.80 30.15 7.75 ;
        RECT  28.35 7.25 30.15 7.75 ;
        RECT  29.65 5.40 30.55 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  31.05 2.65 31.75 3.35 ;
        RECT  31.25 2.65 31.75 9.75 ;
        RECT  31.05 8.15 31.75 9.75 ;
        RECT  31.05 5.40 31.95 6.30 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  6.50 8.10 7.20 11.00 ;
        RECT  10.75 8.85 11.45 11.00 ;
        RECT  16.80 8.20 17.50 11.00 ;
        RECT  19.30 9.55 20.00 11.00 ;
        RECT  24.15 9.30 24.85 11.00 ;
        RECT  26.85 9.30 27.55 11.00 ;
        RECT  29.70 8.25 30.40 11.00 ;
        RECT  0.00 11.00 32.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.45 ;
        RECT  6.50 2.00 7.20 4.40 ;
        RECT  10.70 2.00 11.40 3.95 ;
        RECT  15.80 2.00 16.30 4.25 ;
        RECT  16.90 3.75 17.60 4.95 ;
        RECT  15.80 3.75 20.60 4.25 ;
        RECT  19.90 3.75 20.60 5.45 ;
        RECT  25.55 3.75 26.25 5.45 ;
        RECT  24.60 4.70 26.25 5.45 ;
        RECT  27.35 2.00 27.85 4.25 ;
        RECT  25.55 3.75 27.85 4.25 ;
        RECT  29.70 2.00 30.40 3.30 ;
        RECT  0.00 0.00 32.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.15 3.95 5.20 4.45 ;
        RECT  23.95 6.05 29.15 6.50 ;
        RECT  0.45 3.75 0.95 9.90 ;
        RECT  0.45 3.75 1.15 4.45 ;
        RECT  0.45 8.10 1.15 9.90 ;
        RECT  3.50 6.85 4.20 7.55 ;
        RECT  0.45 7.05 4.20 7.55 ;
        RECT  4.70 3.75 4.85 9.90 ;
        RECT  4.15 8.15 4.85 9.90 ;
        RECT  4.70 3.75 5.05 8.65 ;
        RECT  4.15 3.75 5.05 4.45 ;
        RECT  4.70 3.95 5.20 8.65 ;
        RECT  4.15 8.15 5.20 8.65 ;
        RECT  7.85 3.80 8.55 4.95 ;
        RECT  7.85 7.70 8.55 9.85 ;
        RECT  7.85 4.45 9.30 4.95 ;
        RECT  7.85 7.70 9.25 8.40 ;
        RECT  8.60 4.45 9.30 5.55 ;
        RECT  9.35 3.25 10.25 3.95 ;
        RECT  9.45 6.40 10.15 7.25 ;
        RECT  4.70 6.75 10.15 7.25 ;
        RECT  9.75 3.25 10.25 5.20 ;
        RECT  9.80 7.90 10.30 9.85 ;
        RECT  9.35 9.15 10.30 9.85 ;
        RECT  9.75 4.70 11.10 5.20 ;
        RECT  10.60 4.70 11.10 8.40 ;
        RECT  9.80 7.90 11.10 8.40 ;
        RECT  10.60 6.05 13.15 6.55 ;
        RECT  12.45 6.05 13.15 6.75 ;
        RECT  13.45 4.80 14.15 5.50 ;
        RECT  13.65 4.80 14.15 7.55 ;
        RECT  13.65 6.85 14.40 7.55 ;
        RECT  13.10 3.20 15.35 3.90 ;
        RECT  14.85 3.20 15.35 9.40 ;
        RECT  13.25 8.70 15.35 9.40 ;
        RECT  16.35 5.65 17.05 6.35 ;
        RECT  17.35 6.90 18.05 7.60 ;
        RECT  14.85 7.10 18.05 7.60 ;
        RECT  18.40 4.75 19.10 6.15 ;
        RECT  16.35 5.65 19.10 6.15 ;
        RECT  18.60 4.75 19.10 8.85 ;
        RECT  18.15 8.10 19.10 8.85 ;
        RECT  22.25 4.75 22.50 10.05 ;
        RECT  21.80 7.30 22.50 10.05 ;
        RECT  22.25 4.75 22.75 7.80 ;
        RECT  22.25 4.75 22.95 5.45 ;
        RECT  23.95 6.00 24.65 6.70 ;
        RECT  25.50 8.30 26.20 9.95 ;
        RECT  26.15 7.10 26.85 7.80 ;
        RECT  21.80 7.30 26.85 7.80 ;
        RECT  27.35 6.00 27.85 8.80 ;
        RECT  25.50 8.30 27.85 8.80 ;
        RECT  27.90 4.80 28.60 6.75 ;
        RECT  23.95 6.00 28.60 6.50 ;
        RECT  27.35 6.05 29.15 6.75 ;
    END
END SDFFSX1
MACRO SDFFSX2
    CLASS CORE ;
    FOREIGN SDFFSX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 32.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  16.75 2.55 23.55 3.25 ;
        RECT  22.65 2.55 23.55 3.75 ;
        RECT  16.75 2.55 26.70 3.05 ;
        RECT  26.00 2.55 26.70 3.25 ;
        END
    END SN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  1.45 5.60 2.55 6.30 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END SD
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  28.35 2.65 29.05 4.30 ;
        RECT  28.35 7.25 29.05 10.35 ;
        RECT  28.35 3.80 30.15 4.30 ;
        RECT  29.65 3.80 30.15 7.75 ;
        RECT  28.35 7.25 30.15 7.75 ;
        RECT  29.65 5.40 30.55 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  31.05 2.65 31.75 3.35 ;
        RECT  31.25 2.65 31.75 10.35 ;
        RECT  31.05 8.10 31.75 10.35 ;
        RECT  31.05 5.40 31.95 6.30 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  6.50 8.10 7.20 11.00 ;
        RECT  10.75 8.85 11.45 11.00 ;
        RECT  16.80 8.20 17.50 11.00 ;
        RECT  19.30 9.55 20.00 11.00 ;
        RECT  24.15 9.30 24.85 11.00 ;
        RECT  26.85 9.30 27.55 11.00 ;
        RECT  29.70 8.25 30.40 11.00 ;
        RECT  0.00 11.00 32.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.45 ;
        RECT  6.50 2.00 7.20 4.40 ;
        RECT  10.70 2.00 11.40 3.95 ;
        RECT  15.80 2.00 16.30 4.25 ;
        RECT  16.90 3.75 17.60 4.95 ;
        RECT  15.80 3.75 20.60 4.25 ;
        RECT  19.90 3.75 20.60 5.45 ;
        RECT  25.55 3.75 26.25 5.45 ;
        RECT  24.60 4.70 26.25 5.45 ;
        RECT  27.35 2.00 27.85 4.25 ;
        RECT  25.55 3.75 27.85 4.25 ;
        RECT  29.70 2.00 30.40 3.30 ;
        RECT  0.00 0.00 32.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.15 3.95 5.20 4.45 ;
        RECT  23.95 6.05 29.15 6.50 ;
        RECT  0.45 3.75 0.95 9.90 ;
        RECT  0.45 3.75 1.15 4.45 ;
        RECT  0.45 8.10 1.15 9.90 ;
        RECT  3.50 6.85 4.20 7.55 ;
        RECT  0.45 7.05 4.20 7.55 ;
        RECT  4.70 3.75 4.85 9.90 ;
        RECT  4.15 8.15 4.85 9.90 ;
        RECT  4.70 3.75 5.05 8.65 ;
        RECT  4.15 3.75 5.05 4.45 ;
        RECT  4.70 3.95 5.20 8.65 ;
        RECT  4.15 8.15 5.20 8.65 ;
        RECT  7.85 3.80 8.55 4.95 ;
        RECT  7.85 7.70 8.55 9.85 ;
        RECT  7.85 4.45 9.30 4.95 ;
        RECT  7.85 7.70 9.25 8.40 ;
        RECT  8.60 4.45 9.30 5.55 ;
        RECT  9.35 3.25 10.25 3.95 ;
        RECT  9.45 6.40 10.15 7.25 ;
        RECT  4.70 6.75 10.15 7.25 ;
        RECT  9.75 3.25 10.25 5.20 ;
        RECT  9.80 7.90 10.30 9.85 ;
        RECT  9.35 9.15 10.30 9.85 ;
        RECT  9.75 4.70 11.10 5.20 ;
        RECT  10.60 4.70 11.10 8.40 ;
        RECT  9.80 7.90 11.10 8.40 ;
        RECT  10.60 6.05 13.15 6.55 ;
        RECT  12.45 6.05 13.15 6.75 ;
        RECT  13.45 4.80 14.15 5.50 ;
        RECT  13.65 4.80 14.15 7.55 ;
        RECT  13.65 6.85 14.40 7.55 ;
        RECT  13.10 3.20 15.35 3.90 ;
        RECT  14.85 3.20 15.35 9.40 ;
        RECT  13.25 8.70 15.35 9.40 ;
        RECT  16.35 5.65 17.05 6.35 ;
        RECT  17.35 6.90 18.05 7.60 ;
        RECT  14.85 7.10 18.05 7.60 ;
        RECT  18.40 4.75 19.10 6.15 ;
        RECT  16.35 5.65 19.10 6.15 ;
        RECT  18.60 4.75 19.10 8.85 ;
        RECT  18.15 8.10 19.10 8.85 ;
        RECT  22.25 4.75 22.50 10.05 ;
        RECT  21.80 7.30 22.50 10.05 ;
        RECT  22.25 4.75 22.75 7.80 ;
        RECT  22.25 4.75 22.95 5.45 ;
        RECT  23.95 6.00 24.65 6.70 ;
        RECT  25.50 8.30 26.20 9.95 ;
        RECT  26.15 7.10 26.85 7.80 ;
        RECT  21.80 7.30 26.85 7.80 ;
        RECT  27.35 6.00 27.85 8.80 ;
        RECT  25.50 8.30 27.85 8.80 ;
        RECT  27.90 4.80 28.60 6.75 ;
        RECT  23.95 6.00 28.60 6.50 ;
        RECT  27.35 6.05 29.15 6.75 ;
    END
END SDFFSX2
MACRO SDFFSX4
    CLASS CORE ;
    FOREIGN SDFFSX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 35.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  16.75 2.55 23.55 3.25 ;
        RECT  22.65 2.55 23.55 3.75 ;
        RECT  16.75 2.55 26.70 3.05 ;
        RECT  26.00 2.55 26.70 3.25 ;
        END
    END SN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  1.45 5.60 2.55 6.30 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END SD
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  29.80 2.50 30.30 10.50 ;
        RECT  29.80 2.50 30.50 4.10 ;
        RECT  29.80 8.10 30.50 10.50 ;
        RECT  29.65 5.35 30.55 6.35 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  32.50 2.50 33.20 4.10 ;
        RECT  32.70 2.50 33.20 10.50 ;
        RECT  32.50 5.35 33.20 10.50 ;
        RECT  32.35 5.35 33.35 6.35 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  6.50 8.10 7.20 11.00 ;
        RECT  10.75 8.85 11.45 11.00 ;
        RECT  16.80 8.20 17.50 11.00 ;
        RECT  19.30 9.55 20.00 11.00 ;
        RECT  24.15 9.30 24.85 11.00 ;
        RECT  26.85 9.30 27.55 11.00 ;
        RECT  28.45 8.10 29.15 11.00 ;
        RECT  31.15 8.10 31.85 11.00 ;
        RECT  33.85 8.10 34.55 11.00 ;
        RECT  0.00 11.00 35.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.45 ;
        RECT  6.50 2.00 7.20 4.40 ;
        RECT  10.70 2.00 11.40 3.95 ;
        RECT  15.80 2.00 16.30 4.25 ;
        RECT  16.90 3.75 17.60 4.95 ;
        RECT  15.80 3.75 20.60 4.25 ;
        RECT  19.90 3.75 20.60 5.45 ;
        RECT  25.55 3.75 26.25 5.45 ;
        RECT  24.60 4.70 26.25 5.45 ;
        RECT  28.30 2.00 29.00 4.25 ;
        RECT  25.55 3.75 29.00 4.25 ;
        RECT  31.15 2.00 31.85 4.10 ;
        RECT  33.85 2.00 34.55 4.10 ;
        RECT  0.00 0.00 35.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.15 3.95 5.20 4.45 ;
        RECT  23.95 6.05 29.15 6.50 ;
        RECT  0.45 3.75 0.95 9.90 ;
        RECT  0.45 3.75 1.15 4.45 ;
        RECT  0.45 8.10 1.15 9.90 ;
        RECT  3.50 6.85 4.20 7.55 ;
        RECT  0.45 7.05 4.20 7.55 ;
        RECT  4.70 3.75 4.85 9.90 ;
        RECT  4.15 8.15 4.85 9.90 ;
        RECT  4.70 3.75 5.05 8.65 ;
        RECT  4.15 3.75 5.05 4.45 ;
        RECT  4.70 3.95 5.20 8.65 ;
        RECT  4.15 8.15 5.20 8.65 ;
        RECT  7.85 3.80 8.55 4.95 ;
        RECT  7.85 7.70 8.55 9.85 ;
        RECT  7.85 4.45 9.30 4.95 ;
        RECT  7.85 7.70 9.25 8.40 ;
        RECT  8.60 4.45 9.30 5.55 ;
        RECT  9.35 3.25 10.25 3.95 ;
        RECT  9.45 6.40 10.15 7.25 ;
        RECT  4.70 6.75 10.15 7.25 ;
        RECT  9.75 3.25 10.25 5.20 ;
        RECT  9.80 7.90 10.30 9.85 ;
        RECT  9.35 9.15 10.30 9.85 ;
        RECT  9.75 4.70 11.10 5.20 ;
        RECT  10.60 4.70 11.10 8.40 ;
        RECT  9.80 7.90 11.10 8.40 ;
        RECT  10.60 6.05 13.15 6.55 ;
        RECT  12.45 6.05 13.15 6.75 ;
        RECT  13.45 4.80 14.15 5.50 ;
        RECT  13.65 4.80 14.15 7.55 ;
        RECT  13.65 6.85 14.40 7.55 ;
        RECT  13.10 3.20 15.35 3.90 ;
        RECT  14.85 3.20 15.35 9.40 ;
        RECT  13.25 8.70 15.35 9.40 ;
        RECT  16.35 5.65 17.05 6.35 ;
        RECT  17.35 6.90 18.05 7.60 ;
        RECT  14.85 7.10 18.05 7.60 ;
        RECT  18.40 4.75 19.10 6.15 ;
        RECT  16.35 5.65 19.10 6.15 ;
        RECT  18.60 4.75 19.10 8.85 ;
        RECT  18.15 8.10 19.10 8.85 ;
        RECT  22.25 4.75 22.50 10.05 ;
        RECT  21.80 7.30 22.50 10.05 ;
        RECT  22.25 4.75 22.75 7.80 ;
        RECT  22.25 4.75 22.95 5.45 ;
        RECT  23.95 6.00 24.65 6.70 ;
        RECT  25.50 8.30 26.20 9.95 ;
        RECT  26.15 7.10 26.85 7.80 ;
        RECT  21.80 7.30 26.85 7.80 ;
        RECT  27.35 6.00 27.85 8.80 ;
        RECT  25.50 8.30 27.85 8.80 ;
        RECT  27.90 4.80 28.60 6.75 ;
        RECT  23.95 6.00 28.60 6.50 ;
        RECT  27.35 6.05 29.15 6.75 ;
    END
END SDFFSX4
MACRO SDFFX1
    CLASS CORE ;
    FOREIGN SDFFX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 28.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  1.45 5.60 2.55 6.30 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END SD
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  26.85 3.75 27.55 4.45 ;
        RECT  27.05 3.75 27.55 8.85 ;
        RECT  26.85 7.15 27.55 8.85 ;
        RECT  26.85 5.40 27.75 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  24.15 3.75 24.85 4.45 ;
        RECT  24.30 3.75 24.85 8.85 ;
        RECT  24.15 7.15 24.85 8.85 ;
        RECT  24.05 5.40 24.95 6.30 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  21.45 8.60 22.30 9.10 ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  6.50 8.10 7.20 11.00 ;
        RECT  10.75 8.85 11.45 11.00 ;
        RECT  15.55 8.35 16.25 11.00 ;
        RECT  15.45 9.45 16.25 11.00 ;
        RECT  17.95 10.40 18.65 11.00 ;
        RECT  21.25 7.40 21.95 8.15 ;
        RECT  21.80 7.40 21.95 11.00 ;
        RECT  21.45 7.40 21.95 9.10 ;
        RECT  21.80 8.60 22.30 11.00 ;
        RECT  21.80 10.15 23.50 11.00 ;
        RECT  25.50 7.15 26.20 11.00 ;
        RECT  24.30 10.70 27.55 11.00 ;
        RECT  0.00 11.00 28.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.45 ;
        RECT  6.50 2.00 7.20 4.40 ;
        RECT  10.70 2.00 11.40 3.95 ;
        RECT  15.75 2.00 16.45 4.90 ;
        RECT  21.25 2.00 21.95 3.95 ;
        RECT  25.50 2.00 26.20 4.45 ;
        RECT  0.00 0.00 28.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.15 3.95 5.20 4.45 ;
        RECT  0.45 3.75 0.95 9.90 ;
        RECT  0.45 3.75 1.15 4.45 ;
        RECT  0.45 8.10 1.15 9.90 ;
        RECT  3.50 6.85 4.20 7.55 ;
        RECT  0.45 7.05 4.20 7.55 ;
        RECT  4.70 3.75 4.85 9.90 ;
        RECT  4.15 8.15 4.85 9.90 ;
        RECT  4.70 3.75 5.05 8.65 ;
        RECT  4.15 3.75 5.05 4.45 ;
        RECT  4.70 3.95 5.20 8.65 ;
        RECT  4.15 8.15 5.20 8.65 ;
        RECT  7.85 3.80 8.55 4.95 ;
        RECT  7.85 7.70 8.55 9.85 ;
        RECT  7.85 4.45 9.30 4.95 ;
        RECT  7.85 7.70 9.25 8.40 ;
        RECT  8.60 4.45 9.30 5.55 ;
        RECT  9.35 3.25 10.25 3.95 ;
        RECT  9.45 6.40 10.15 7.25 ;
        RECT  4.70 6.75 10.15 7.25 ;
        RECT  9.75 3.25 10.25 5.20 ;
        RECT  9.80 7.90 10.30 9.85 ;
        RECT  9.35 9.15 10.30 9.85 ;
        RECT  9.75 4.70 11.10 5.20 ;
        RECT  10.60 4.70 11.10 8.40 ;
        RECT  9.80 7.90 11.10 8.40 ;
        RECT  10.60 6.05 13.15 6.55 ;
        RECT  12.45 6.05 13.15 6.75 ;
        RECT  12.65 7.30 13.35 8.00 ;
        RECT  13.45 4.80 14.15 5.50 ;
        RECT  13.10 8.45 13.80 10.15 ;
        RECT  13.65 4.80 14.15 7.80 ;
        RECT  12.65 7.30 14.15 7.80 ;
        RECT  13.10 3.25 15.10 3.95 ;
        RECT  14.60 3.25 15.10 8.95 ;
        RECT  13.10 8.45 15.10 8.95 ;
        RECT  15.55 5.45 16.25 6.15 ;
        RECT  14.60 6.70 17.00 7.20 ;
        RECT  16.30 6.70 17.00 7.40 ;
        RECT  17.25 4.15 17.95 4.85 ;
        RECT  15.55 5.45 17.95 5.95 ;
        RECT  17.45 4.15 17.95 9.05 ;
        RECT  16.95 8.35 17.95 9.05 ;
        RECT  18.90 3.30 19.60 4.00 ;
        RECT  19.10 3.30 19.60 10.15 ;
        RECT  19.10 9.65 21.00 10.15 ;
        RECT  20.30 9.65 21.00 10.35 ;
        RECT  20.80 4.45 21.50 5.15 ;
        RECT  21.60 5.70 22.30 6.40 ;
        RECT  19.10 5.90 22.30 6.40 ;
        RECT  22.60 3.25 23.30 3.95 ;
        RECT  20.80 4.45 23.30 4.95 ;
        RECT  22.60 7.40 23.30 8.15 ;
        RECT  22.80 3.25 23.30 9.65 ;
        RECT  22.80 8.95 23.65 9.65 ;
    END
END SDFFX1
MACRO SDFFX2
    CLASS CORE ;
    FOREIGN SDFFX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 28.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  1.45 5.60 2.55 6.30 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END SD
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  26.85 2.70 27.55 4.50 ;
        RECT  27.05 2.70 27.55 10.55 ;
        RECT  26.85 7.10 27.55 10.55 ;
        RECT  26.85 5.40 27.75 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  24.15 2.70 24.85 4.50 ;
        RECT  24.30 2.70 24.85 10.55 ;
        RECT  24.15 7.10 24.85 10.55 ;
        RECT  24.05 5.40 24.95 6.30 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  6.50 8.10 7.20 11.00 ;
        RECT  10.75 8.85 11.45 11.00 ;
        RECT  15.55 8.35 16.25 11.00 ;
        RECT  15.45 9.45 16.25 11.00 ;
        RECT  17.95 10.40 18.65 11.00 ;
        RECT  21.25 7.40 21.95 8.15 ;
        RECT  21.45 7.40 21.95 11.00 ;
        RECT  25.50 7.10 26.20 11.00 ;
        RECT  0.00 11.00 28.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.45 ;
        RECT  6.50 2.00 7.20 4.40 ;
        RECT  10.70 2.00 11.40 3.95 ;
        RECT  15.75 2.00 16.45 4.90 ;
        RECT  21.25 2.00 21.95 3.95 ;
        RECT  25.50 2.00 26.20 4.50 ;
        RECT  0.00 0.00 28.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.15 3.95 5.20 4.45 ;
        RECT  0.45 3.75 0.95 9.90 ;
        RECT  0.45 3.75 1.15 4.45 ;
        RECT  0.45 8.10 1.15 9.90 ;
        RECT  3.50 6.85 4.20 7.55 ;
        RECT  0.45 7.05 4.20 7.55 ;
        RECT  4.70 3.75 4.85 9.90 ;
        RECT  4.15 8.15 4.85 9.90 ;
        RECT  4.70 3.75 5.05 8.65 ;
        RECT  4.15 3.75 5.05 4.45 ;
        RECT  4.70 3.95 5.20 8.65 ;
        RECT  4.15 8.15 5.20 8.65 ;
        RECT  7.85 3.80 8.55 4.95 ;
        RECT  7.85 7.70 8.55 9.85 ;
        RECT  7.85 4.45 9.30 4.95 ;
        RECT  7.85 7.70 9.25 8.40 ;
        RECT  8.60 4.45 9.30 5.55 ;
        RECT  9.35 3.25 10.25 3.95 ;
        RECT  9.45 6.40 10.15 7.25 ;
        RECT  4.70 6.75 10.15 7.25 ;
        RECT  9.75 3.25 10.25 5.20 ;
        RECT  9.80 7.90 10.30 9.85 ;
        RECT  9.35 9.15 10.30 9.85 ;
        RECT  9.75 4.70 11.10 5.20 ;
        RECT  10.60 4.70 11.10 8.40 ;
        RECT  9.80 7.90 11.10 8.40 ;
        RECT  10.60 6.05 13.15 6.55 ;
        RECT  12.45 6.05 13.15 6.75 ;
        RECT  12.65 7.30 13.35 8.00 ;
        RECT  13.45 4.80 14.15 5.50 ;
        RECT  13.10 8.45 13.80 10.15 ;
        RECT  13.65 4.80 14.15 7.80 ;
        RECT  12.65 7.30 14.15 7.80 ;
        RECT  13.10 3.25 15.10 3.95 ;
        RECT  14.60 3.25 15.10 8.95 ;
        RECT  13.10 8.45 15.10 8.95 ;
        RECT  15.55 5.45 16.25 6.15 ;
        RECT  14.60 6.70 17.00 7.20 ;
        RECT  16.30 6.70 17.00 7.40 ;
        RECT  17.25 4.15 17.95 4.85 ;
        RECT  15.55 5.45 17.95 5.95 ;
        RECT  17.45 4.15 17.95 9.05 ;
        RECT  16.95 8.35 17.95 9.05 ;
        RECT  18.90 3.30 19.60 4.00 ;
        RECT  19.10 3.30 19.60 10.15 ;
        RECT  19.10 9.65 21.00 10.15 ;
        RECT  20.30 9.65 21.00 10.35 ;
        RECT  20.80 4.45 21.50 5.15 ;
        RECT  21.60 5.70 22.30 6.40 ;
        RECT  19.10 5.90 22.30 6.40 ;
        RECT  22.60 3.25 23.30 3.95 ;
        RECT  20.80 4.45 23.30 4.95 ;
        RECT  22.60 7.40 23.30 8.15 ;
        RECT  22.80 3.25 23.30 9.65 ;
        RECT  22.80 8.95 23.65 9.65 ;
    END
END SDFFX2
MACRO SDFFX4
    CLASS CORE ;
    FOREIGN SDFFX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 30.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  1.45 5.60 2.55 6.30 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END SD
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  28.30 2.90 29.00 4.50 ;
        RECT  28.50 2.90 29.00 10.50 ;
        RECT  28.30 5.35 29.00 10.50 ;
        RECT  28.15 5.35 29.15 6.35 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  25.60 2.90 26.10 10.50 ;
        RECT  25.60 2.90 26.30 4.50 ;
        RECT  25.60 7.10 26.30 10.50 ;
        RECT  25.45 5.35 26.35 6.35 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  6.50 8.10 7.20 11.00 ;
        RECT  10.75 8.85 11.45 11.00 ;
        RECT  15.55 8.35 16.25 11.00 ;
        RECT  15.45 9.45 16.25 11.00 ;
        RECT  17.95 10.40 18.65 11.00 ;
        RECT  21.25 7.40 21.95 8.15 ;
        RECT  21.45 7.40 21.95 11.00 ;
        RECT  24.25 7.10 24.95 11.00 ;
        RECT  26.95 7.10 27.65 11.00 ;
        RECT  29.65 7.10 30.35 11.00 ;
        RECT  0.00 11.00 30.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.45 ;
        RECT  6.50 2.00 7.20 4.40 ;
        RECT  10.70 2.00 11.40 3.95 ;
        RECT  15.75 2.00 16.45 4.90 ;
        RECT  21.25 2.00 21.95 3.95 ;
        RECT  24.25 2.00 24.95 4.50 ;
        RECT  26.95 2.00 27.65 4.50 ;
        RECT  29.65 2.00 30.35 4.50 ;
        RECT  0.00 0.00 30.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.15 3.95 5.20 4.45 ;
        RECT  0.45 3.75 0.95 9.90 ;
        RECT  0.45 3.75 1.15 4.45 ;
        RECT  0.45 8.10 1.15 9.90 ;
        RECT  3.50 6.85 4.20 7.55 ;
        RECT  0.45 7.05 4.20 7.55 ;
        RECT  4.70 3.75 4.85 9.90 ;
        RECT  4.15 8.15 4.85 9.90 ;
        RECT  4.70 3.75 5.05 8.65 ;
        RECT  4.15 3.75 5.05 4.45 ;
        RECT  4.70 3.95 5.20 8.65 ;
        RECT  4.15 8.15 5.20 8.65 ;
        RECT  7.85 3.80 8.55 4.95 ;
        RECT  7.85 7.70 8.55 9.85 ;
        RECT  7.85 4.45 9.30 4.95 ;
        RECT  7.85 7.70 9.25 8.40 ;
        RECT  8.60 4.45 9.30 5.55 ;
        RECT  9.35 3.25 10.25 3.95 ;
        RECT  9.45 6.40 10.15 7.25 ;
        RECT  4.70 6.75 10.15 7.25 ;
        RECT  9.75 3.25 10.25 5.20 ;
        RECT  9.80 7.90 10.30 9.85 ;
        RECT  9.35 9.15 10.30 9.85 ;
        RECT  9.75 4.70 11.10 5.20 ;
        RECT  10.60 4.70 11.10 8.40 ;
        RECT  9.80 7.90 11.10 8.40 ;
        RECT  10.60 6.05 13.15 6.55 ;
        RECT  12.45 6.05 13.15 6.75 ;
        RECT  12.65 7.30 13.35 8.00 ;
        RECT  13.45 4.80 14.15 5.50 ;
        RECT  13.10 8.45 13.80 10.15 ;
        RECT  13.65 4.80 14.15 7.80 ;
        RECT  12.65 7.30 14.15 7.80 ;
        RECT  13.10 3.25 15.10 3.95 ;
        RECT  14.60 3.25 15.10 8.95 ;
        RECT  13.10 8.45 15.10 8.95 ;
        RECT  15.55 5.45 16.25 6.15 ;
        RECT  14.60 6.70 17.00 7.20 ;
        RECT  16.30 6.70 17.00 7.40 ;
        RECT  17.25 4.15 17.95 4.85 ;
        RECT  15.55 5.45 17.95 5.95 ;
        RECT  17.45 4.15 17.95 9.05 ;
        RECT  16.95 8.35 17.95 9.05 ;
        RECT  18.90 3.30 19.60 4.00 ;
        RECT  19.10 3.30 19.60 10.15 ;
        RECT  19.10 9.65 21.00 10.15 ;
        RECT  20.30 9.65 21.00 10.35 ;
        RECT  20.80 4.45 21.50 5.15 ;
        RECT  21.60 5.70 22.30 6.40 ;
        RECT  19.10 5.90 22.30 6.40 ;
        RECT  22.60 3.25 23.30 3.95 ;
        RECT  20.80 4.45 23.30 4.95 ;
        RECT  22.60 7.40 23.30 8.15 ;
        RECT  22.80 3.25 23.30 9.65 ;
        RECT  22.80 8.95 23.65 9.65 ;
    END
END SDFFX4
MACRO SDFRRSX1
    CLASS CORE ;
    FOREIGN SDFRRSX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 35.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  16.50 2.55 17.95 3.25 ;
        RECT  17.05 2.55 17.95 3.75 ;
        RECT  16.50 2.55 29.50 3.05 ;
        RECT  28.80 2.55 29.50 3.25 ;
        END
    END SN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  1.45 5.60 2.55 6.30 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END SD
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  20.45 5.75 21.15 6.45 ;
        RECT  22.65 5.35 23.55 6.35 ;
        RECT  20.45 5.85 23.55 6.35 ;
        RECT  22.65 5.50 24.90 6.20 ;
        RECT  20.45 5.85 24.90 6.20 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  31.15 2.65 31.85 4.30 ;
        RECT  31.15 7.25 31.85 9.75 ;
        RECT  31.15 3.80 32.95 4.30 ;
        RECT  32.45 3.80 32.95 7.75 ;
        RECT  31.15 7.25 32.95 7.75 ;
        RECT  32.45 5.35 33.35 6.35 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  33.85 2.65 34.55 3.35 ;
        RECT  34.05 2.65 34.55 9.75 ;
        RECT  33.85 7.95 34.55 9.75 ;
        RECT  33.75 7.95 34.75 8.95 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  6.50 8.10 7.20 11.00 ;
        RECT  11.05 9.00 11.75 11.00 ;
        RECT  16.80 8.45 17.50 11.00 ;
        RECT  19.65 7.30 20.35 11.00 ;
        RECT  19.65 7.30 25.35 7.80 ;
        RECT  24.65 7.30 25.35 8.35 ;
        RECT  26.85 9.25 27.55 11.00 ;
        RECT  29.55 9.25 30.25 11.00 ;
        RECT  32.50 8.25 33.20 11.00 ;
        RECT  0.00 11.00 35.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.45 ;
        RECT  6.50 2.00 7.20 4.40 ;
        RECT  11.05 2.00 11.75 4.85 ;
        RECT  15.50 2.00 16.00 4.80 ;
        RECT  16.90 4.30 17.60 5.05 ;
        RECT  18.45 3.55 18.95 4.80 ;
        RECT  15.50 4.30 18.95 4.80 ;
        RECT  18.45 3.55 21.85 4.05 ;
        RECT  21.15 3.55 21.85 4.25 ;
        RECT  26.85 3.55 27.55 4.25 ;
        RECT  26.85 3.75 30.65 4.25 ;
        RECT  30.15 2.00 30.65 5.50 ;
        RECT  30.15 4.80 31.40 5.50 ;
        RECT  32.50 2.00 33.20 3.30 ;
        RECT  0.00 0.00 35.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.15 3.95 5.20 4.45 ;
        RECT  7.85 9.60 9.70 9.95 ;
        RECT  0.45 3.75 0.95 9.90 ;
        RECT  0.45 3.75 1.15 4.45 ;
        RECT  0.45 8.10 1.15 9.90 ;
        RECT  3.50 6.85 4.20 7.55 ;
        RECT  0.45 7.05 4.20 7.55 ;
        RECT  4.70 3.75 4.85 9.90 ;
        RECT  4.15 8.15 4.85 9.90 ;
        RECT  4.70 3.75 5.05 8.65 ;
        RECT  4.15 3.75 5.05 4.45 ;
        RECT  4.70 3.95 5.20 8.65 ;
        RECT  4.15 8.15 5.20 8.65 ;
        RECT  8.15 8.10 8.55 10.30 ;
        RECT  7.85 8.10 8.55 9.95 ;
        RECT  7.85 3.75 9.20 4.50 ;
        RECT  8.70 3.75 9.20 6.35 ;
        RECT  8.70 5.65 9.55 6.35 ;
        RECT  8.15 9.60 9.70 10.30 ;
        RECT  9.70 4.20 10.55 4.90 ;
        RECT  9.70 8.00 10.40 9.00 ;
        RECT  10.05 4.20 10.55 6.05 ;
        RECT  11.50 6.65 12.20 7.35 ;
        RECT  4.70 6.85 12.20 7.35 ;
        RECT  10.05 5.55 13.35 6.05 ;
        RECT  12.35 3.20 12.85 6.05 ;
        RECT  12.85 5.55 13.35 8.50 ;
        RECT  9.70 8.00 13.35 8.50 ;
        RECT  12.85 6.70 13.55 7.40 ;
        RECT  13.40 4.20 14.55 4.90 ;
        RECT  13.85 3.00 14.55 3.70 ;
        RECT  12.35 3.20 14.55 3.70 ;
        RECT  14.05 4.20 14.55 9.70 ;
        RECT  13.40 9.00 15.00 9.70 ;
        RECT  16.35 5.65 17.05 6.35 ;
        RECT  17.35 7.25 18.05 7.95 ;
        RECT  14.05 7.45 18.05 7.95 ;
        RECT  18.65 5.65 19.15 9.15 ;
        RECT  18.15 8.45 19.15 9.15 ;
        RECT  19.45 4.55 19.95 6.15 ;
        RECT  16.35 5.65 19.95 6.15 ;
        RECT  19.45 4.55 20.15 5.25 ;
        RECT  22.00 8.30 22.70 10.05 ;
        RECT  23.50 3.55 24.20 4.25 ;
        RECT  24.50 8.85 25.20 9.95 ;
        RECT  23.50 3.75 26.35 4.25 ;
        RECT  25.85 3.75 26.35 9.35 ;
        RECT  22.00 8.85 26.35 9.35 ;
        RECT  26.85 4.75 29.05 5.45 ;
        RECT  28.20 8.25 28.90 9.90 ;
        RECT  28.55 4.75 29.05 6.55 ;
        RECT  28.95 7.05 29.65 7.75 ;
        RECT  25.85 7.25 29.65 7.75 ;
        RECT  30.15 6.05 30.65 8.75 ;
        RECT  28.20 8.25 30.65 8.75 ;
        RECT  28.55 6.05 31.95 6.55 ;
        RECT  31.25 6.05 31.95 6.75 ;
    END
END SDFRRSX1
MACRO SDFRRSX2
    CLASS CORE ;
    FOREIGN SDFRRSX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 35.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  16.50 2.55 17.95 3.25 ;
        RECT  17.05 2.55 17.95 3.75 ;
        RECT  16.50 2.55 29.50 3.05 ;
        RECT  28.80 2.55 29.50 3.25 ;
        END
    END SN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  1.45 5.60 2.55 6.30 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END SD
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  20.45 5.75 21.15 6.45 ;
        RECT  22.65 5.35 23.55 6.35 ;
        RECT  20.45 5.85 23.55 6.35 ;
        RECT  22.65 5.50 24.90 6.20 ;
        RECT  20.45 5.85 24.90 6.20 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  31.15 2.65 31.85 4.30 ;
        RECT  31.15 7.25 31.85 10.50 ;
        RECT  31.15 3.80 32.95 4.30 ;
        RECT  32.45 3.80 32.95 7.75 ;
        RECT  31.15 7.25 32.95 7.75 ;
        RECT  32.45 5.35 33.35 6.35 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  33.85 2.65 34.55 3.35 ;
        RECT  34.05 2.65 34.55 10.50 ;
        RECT  33.85 7.95 34.55 10.50 ;
        RECT  33.75 7.95 34.75 8.95 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  6.50 8.10 7.20 11.00 ;
        RECT  11.05 9.00 11.75 11.00 ;
        RECT  16.80 8.45 17.50 11.00 ;
        RECT  19.65 7.30 20.35 11.00 ;
        RECT  19.65 7.30 25.35 7.80 ;
        RECT  24.65 7.30 25.35 8.35 ;
        RECT  26.85 9.25 27.55 11.00 ;
        RECT  29.55 9.25 30.25 11.00 ;
        RECT  32.50 8.25 33.20 11.00 ;
        RECT  0.00 11.00 35.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.45 ;
        RECT  6.50 2.00 7.20 4.40 ;
        RECT  11.05 2.00 11.75 4.85 ;
        RECT  15.50 2.00 16.00 4.80 ;
        RECT  16.90 4.30 17.60 5.05 ;
        RECT  18.45 3.55 18.95 4.80 ;
        RECT  15.50 4.30 18.95 4.80 ;
        RECT  18.45 3.55 21.85 4.05 ;
        RECT  21.15 3.55 21.85 4.25 ;
        RECT  26.85 3.55 27.55 4.25 ;
        RECT  26.85 3.75 30.65 4.25 ;
        RECT  30.15 2.00 30.65 5.50 ;
        RECT  30.15 4.80 31.40 5.50 ;
        RECT  32.50 2.00 33.20 3.30 ;
        RECT  0.00 0.00 35.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.15 3.95 5.20 4.45 ;
        RECT  7.85 9.60 9.70 9.95 ;
        RECT  0.45 3.75 0.95 9.90 ;
        RECT  0.45 3.75 1.15 4.45 ;
        RECT  0.45 8.10 1.15 9.90 ;
        RECT  3.50 6.85 4.20 7.55 ;
        RECT  0.45 7.05 4.20 7.55 ;
        RECT  4.70 3.75 4.85 9.90 ;
        RECT  4.15 8.15 4.85 9.90 ;
        RECT  4.70 3.75 5.05 8.65 ;
        RECT  4.15 3.75 5.05 4.45 ;
        RECT  4.70 3.95 5.20 8.65 ;
        RECT  4.15 8.15 5.20 8.65 ;
        RECT  8.15 8.10 8.55 10.30 ;
        RECT  7.85 8.10 8.55 9.95 ;
        RECT  7.85 3.75 9.20 4.50 ;
        RECT  8.70 3.75 9.20 6.35 ;
        RECT  8.70 5.65 9.55 6.35 ;
        RECT  8.15 9.60 9.70 10.30 ;
        RECT  9.70 4.20 10.55 4.90 ;
        RECT  9.70 8.00 10.40 9.00 ;
        RECT  10.05 4.20 10.55 6.05 ;
        RECT  11.50 6.65 12.20 7.35 ;
        RECT  4.70 6.85 12.20 7.35 ;
        RECT  10.05 5.55 13.35 6.05 ;
        RECT  12.35 3.20 12.85 6.05 ;
        RECT  12.85 5.55 13.35 8.50 ;
        RECT  9.70 8.00 13.35 8.50 ;
        RECT  12.85 6.70 13.55 7.40 ;
        RECT  13.40 4.20 14.55 4.90 ;
        RECT  13.85 3.00 14.55 3.70 ;
        RECT  12.35 3.20 14.55 3.70 ;
        RECT  14.05 4.20 14.55 9.70 ;
        RECT  13.40 9.00 15.00 9.70 ;
        RECT  16.35 5.65 17.05 6.35 ;
        RECT  17.35 7.25 18.05 7.95 ;
        RECT  14.05 7.45 18.05 7.95 ;
        RECT  18.65 5.65 19.15 9.15 ;
        RECT  18.15 8.45 19.15 9.15 ;
        RECT  19.45 4.55 19.95 6.15 ;
        RECT  16.35 5.65 19.95 6.15 ;
        RECT  19.45 4.55 20.15 5.25 ;
        RECT  22.00 8.30 22.70 10.05 ;
        RECT  23.50 3.55 24.20 4.25 ;
        RECT  24.50 8.85 25.20 9.95 ;
        RECT  23.50 3.75 26.35 4.25 ;
        RECT  25.85 3.75 26.35 9.35 ;
        RECT  22.00 8.85 26.35 9.35 ;
        RECT  26.85 4.75 29.05 5.45 ;
        RECT  28.20 8.25 28.90 9.90 ;
        RECT  28.55 4.75 29.05 6.55 ;
        RECT  28.95 7.05 29.65 7.75 ;
        RECT  25.85 7.25 29.65 7.75 ;
        RECT  30.15 6.05 30.65 8.75 ;
        RECT  28.20 8.25 30.65 8.75 ;
        RECT  28.55 6.05 31.95 6.55 ;
        RECT  31.25 6.05 31.95 6.75 ;
    END
END SDFRRSX2
MACRO SDFRRSX4
    CLASS CORE ;
    FOREIGN SDFRRSX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 37.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  16.50 2.55 17.95 3.25 ;
        RECT  17.05 2.55 17.95 3.75 ;
        RECT  16.50 2.55 29.50 3.05 ;
        RECT  28.80 2.55 29.50 3.25 ;
        END
    END SN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  1.45 5.60 2.55 6.30 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END SD
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  20.45 5.75 21.15 6.45 ;
        RECT  22.65 5.35 23.55 6.35 ;
        RECT  20.45 5.85 23.55 6.35 ;
        RECT  22.65 5.50 24.90 6.20 ;
        RECT  20.45 5.85 24.90 6.20 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  32.60 2.50 33.10 10.50 ;
        RECT  32.60 2.50 33.30 4.10 ;
        RECT  32.60 8.10 33.30 10.50 ;
        RECT  32.45 5.35 33.35 6.35 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  35.30 2.50 36.00 4.10 ;
        RECT  35.50 2.50 36.00 10.50 ;
        RECT  35.30 5.35 36.00 10.50 ;
        RECT  35.15 5.35 36.15 6.35 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  6.50 8.10 7.20 11.00 ;
        RECT  11.05 9.00 11.75 11.00 ;
        RECT  16.80 8.45 17.50 11.00 ;
        RECT  19.65 7.30 20.35 11.00 ;
        RECT  19.65 7.30 25.35 7.80 ;
        RECT  24.65 7.30 25.35 8.35 ;
        RECT  26.85 9.25 27.55 11.00 ;
        RECT  29.55 9.25 30.25 11.00 ;
        RECT  31.25 8.10 31.95 11.00 ;
        RECT  33.95 8.10 34.65 11.00 ;
        RECT  36.65 8.10 37.35 11.00 ;
        RECT  0.00 11.00 37.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.45 ;
        RECT  6.50 2.00 7.20 4.40 ;
        RECT  11.05 2.00 11.75 4.85 ;
        RECT  15.50 2.00 16.00 4.80 ;
        RECT  16.90 4.30 17.60 5.05 ;
        RECT  18.45 3.55 18.95 4.80 ;
        RECT  15.50 4.30 18.95 4.80 ;
        RECT  18.45 3.55 21.85 4.05 ;
        RECT  21.15 3.55 21.85 4.25 ;
        RECT  26.85 3.55 27.55 4.25 ;
        RECT  26.85 3.75 30.60 4.25 ;
        RECT  30.10 2.00 30.60 5.50 ;
        RECT  30.10 4.80 31.40 5.50 ;
        RECT  31.10 2.00 31.80 3.90 ;
        RECT  33.95 2.00 34.65 4.10 ;
        RECT  36.65 2.00 37.35 4.10 ;
        RECT  0.00 0.00 37.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.15 3.95 5.20 4.45 ;
        RECT  7.85 9.60 9.70 9.95 ;
        RECT  0.45 3.75 0.95 9.90 ;
        RECT  0.45 3.75 1.15 4.45 ;
        RECT  0.45 8.10 1.15 9.90 ;
        RECT  3.50 6.85 4.20 7.55 ;
        RECT  0.45 7.05 4.20 7.55 ;
        RECT  4.70 3.75 4.85 9.90 ;
        RECT  4.15 8.15 4.85 9.90 ;
        RECT  4.70 3.75 5.05 8.65 ;
        RECT  4.15 3.75 5.05 4.45 ;
        RECT  4.70 3.95 5.20 8.65 ;
        RECT  4.15 8.15 5.20 8.65 ;
        RECT  8.15 8.10 8.55 10.30 ;
        RECT  7.85 8.10 8.55 9.95 ;
        RECT  7.85 3.75 9.20 4.50 ;
        RECT  8.70 3.75 9.20 6.35 ;
        RECT  8.70 5.65 9.55 6.35 ;
        RECT  8.15 9.60 9.70 10.30 ;
        RECT  9.70 4.20 10.55 4.90 ;
        RECT  9.70 8.00 10.40 9.00 ;
        RECT  10.05 4.20 10.55 6.05 ;
        RECT  11.50 6.65 12.20 7.35 ;
        RECT  4.70 6.85 12.20 7.35 ;
        RECT  10.05 5.55 13.35 6.05 ;
        RECT  12.35 3.20 12.85 6.05 ;
        RECT  12.85 5.55 13.35 8.50 ;
        RECT  9.70 8.00 13.35 8.50 ;
        RECT  12.85 6.70 13.55 7.40 ;
        RECT  13.40 4.20 14.55 4.90 ;
        RECT  13.85 3.00 14.55 3.70 ;
        RECT  12.35 3.20 14.55 3.70 ;
        RECT  14.05 4.20 14.55 9.70 ;
        RECT  13.40 9.00 15.00 9.70 ;
        RECT  16.35 5.65 17.05 6.35 ;
        RECT  17.35 7.25 18.05 7.95 ;
        RECT  14.05 7.45 18.05 7.95 ;
        RECT  18.65 5.65 19.15 9.15 ;
        RECT  18.15 8.45 19.15 9.15 ;
        RECT  19.45 4.55 19.95 6.15 ;
        RECT  16.35 5.65 19.95 6.15 ;
        RECT  19.45 4.55 20.15 5.25 ;
        RECT  22.00 8.30 22.70 10.05 ;
        RECT  23.50 3.55 24.20 4.25 ;
        RECT  24.50 8.85 25.20 9.95 ;
        RECT  23.50 3.75 26.35 4.25 ;
        RECT  25.85 3.75 26.35 9.35 ;
        RECT  22.00 8.85 26.35 9.35 ;
        RECT  26.85 4.75 29.05 5.45 ;
        RECT  28.20 8.25 28.90 9.90 ;
        RECT  28.55 4.75 29.05 6.55 ;
        RECT  28.95 7.05 29.65 7.75 ;
        RECT  25.85 7.25 29.65 7.75 ;
        RECT  30.15 6.05 30.65 8.75 ;
        RECT  28.20 8.25 30.65 8.75 ;
        RECT  28.55 6.05 31.95 6.55 ;
        RECT  31.25 6.05 31.95 6.75 ;
    END
END SDFRRSX4
MACRO SDFRRX1
    CLASS CORE ;
    FOREIGN SDFRRX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 30.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  1.45 5.60 2.55 6.30 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END SD
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  18.45 7.05 19.15 8.40 ;
        RECT  19.85 6.70 20.75 7.60 ;
        RECT  20.25 5.45 20.75 7.60 ;
        RECT  18.45 7.05 20.75 7.60 ;
        RECT  20.90 5.25 21.60 5.95 ;
        RECT  20.25 5.45 21.60 5.95 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  29.65 3.75 30.35 4.45 ;
        RECT  29.85 3.75 30.35 8.85 ;
        RECT  29.65 7.15 30.35 8.85 ;
        RECT  29.65 5.40 30.55 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  26.95 3.75 27.65 4.45 ;
        RECT  27.10 3.75 27.65 8.85 ;
        RECT  26.95 7.15 27.65 8.85 ;
        RECT  26.85 5.40 27.75 6.30 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  6.50 8.10 7.20 11.00 ;
        RECT  11.05 9.00 11.75 11.00 ;
        RECT  15.75 7.90 16.45 11.00 ;
        RECT  19.05 8.90 19.75 11.00 ;
        RECT  24.05 7.40 24.75 11.00 ;
        RECT  28.30 7.15 29.00 11.00 ;
        RECT  24.05 10.70 30.35 11.00 ;
        RECT  0.00 11.00 30.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.45 ;
        RECT  6.50 2.00 7.20 4.40 ;
        RECT  11.05 2.00 11.75 4.85 ;
        RECT  15.15 2.00 16.75 3.15 ;
        RECT  16.05 2.00 16.75 4.90 ;
        RECT  18.20 2.00 18.90 3.25 ;
        RECT  24.05 2.00 24.75 3.95 ;
        RECT  28.30 2.00 29.00 4.45 ;
        RECT  0.00 0.00 30.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.15 3.95 5.20 4.45 ;
        RECT  7.85 9.60 9.70 9.95 ;
        RECT  0.45 3.75 0.95 9.90 ;
        RECT  0.45 3.75 1.15 4.45 ;
        RECT  0.45 8.10 1.15 9.90 ;
        RECT  3.50 6.85 4.20 7.55 ;
        RECT  0.45 7.05 4.20 7.55 ;
        RECT  4.70 3.75 4.85 9.90 ;
        RECT  4.15 8.15 4.85 9.90 ;
        RECT  4.70 3.75 5.05 8.65 ;
        RECT  4.15 3.75 5.05 4.45 ;
        RECT  4.70 3.95 5.20 8.65 ;
        RECT  4.15 8.15 5.20 8.65 ;
        RECT  8.15 8.10 8.55 10.30 ;
        RECT  7.85 8.10 8.55 9.95 ;
        RECT  7.85 3.75 9.20 4.50 ;
        RECT  8.70 3.75 9.20 6.35 ;
        RECT  8.70 5.65 9.55 6.35 ;
        RECT  8.15 9.60 9.70 10.30 ;
        RECT  9.70 4.20 10.55 4.90 ;
        RECT  9.70 8.00 10.40 9.00 ;
        RECT  10.05 4.20 10.55 6.05 ;
        RECT  11.50 6.65 12.20 7.35 ;
        RECT  4.70 6.85 12.20 7.35 ;
        RECT  10.05 5.55 13.35 6.05 ;
        RECT  12.35 3.20 12.85 6.05 ;
        RECT  12.85 5.55 13.35 8.50 ;
        RECT  9.70 8.00 13.35 8.50 ;
        RECT  12.85 6.70 13.55 7.40 ;
        RECT  13.40 4.20 14.10 4.90 ;
        RECT  13.40 4.40 14.55 4.90 ;
        RECT  14.05 4.20 14.10 9.70 ;
        RECT  13.40 9.00 14.10 9.70 ;
        RECT  13.85 3.00 14.55 3.70 ;
        RECT  12.35 3.20 14.55 3.70 ;
        RECT  14.05 4.40 14.55 9.50 ;
        RECT  13.40 9.00 14.55 9.50 ;
        RECT  15.30 5.45 16.00 6.15 ;
        RECT  14.05 6.70 16.95 7.20 ;
        RECT  16.25 6.70 16.95 7.40 ;
        RECT  15.30 5.45 17.95 5.95 ;
        RECT  17.45 4.35 17.95 9.70 ;
        RECT  17.45 9.00 18.25 9.70 ;
        RECT  18.55 4.15 19.25 4.85 ;
        RECT  17.45 4.35 19.25 4.85 ;
        RECT  20.70 3.30 21.40 4.00 ;
        RECT  20.70 3.45 22.60 4.00 ;
        RECT  21.55 7.20 22.10 10.50 ;
        RECT  21.40 8.75 22.10 10.50 ;
        RECT  22.10 3.45 22.60 7.90 ;
        RECT  21.55 7.20 22.60 7.90 ;
        RECT  23.60 4.45 24.30 5.15 ;
        RECT  24.40 5.70 25.10 6.40 ;
        RECT  22.10 5.90 25.10 6.40 ;
        RECT  25.40 3.25 26.10 3.95 ;
        RECT  23.60 4.45 26.10 4.95 ;
        RECT  25.60 3.25 26.10 10.10 ;
        RECT  25.40 7.40 26.10 10.10 ;
    END
END SDFRRX1
MACRO SDFRRX2
    CLASS CORE ;
    FOREIGN SDFRRX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 30.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  1.45 5.60 2.55 6.30 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END SD
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  18.45 7.05 19.15 8.40 ;
        RECT  19.85 6.70 20.75 7.60 ;
        RECT  20.25 5.45 20.75 7.60 ;
        RECT  18.45 7.05 20.75 7.60 ;
        RECT  20.90 5.25 21.60 5.95 ;
        RECT  20.25 5.45 21.60 5.95 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  29.65 2.70 30.35 4.50 ;
        RECT  29.85 2.70 30.35 10.50 ;
        RECT  29.65 7.10 30.35 10.50 ;
        RECT  29.65 5.40 30.55 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  26.95 2.70 27.65 4.50 ;
        RECT  27.10 2.70 27.65 10.50 ;
        RECT  26.95 7.10 27.65 10.50 ;
        RECT  26.85 5.40 27.75 6.30 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  6.50 8.10 7.20 11.00 ;
        RECT  11.05 9.00 11.75 11.00 ;
        RECT  15.75 7.90 16.45 11.00 ;
        RECT  19.05 8.90 19.75 11.00 ;
        RECT  24.05 7.40 24.75 11.00 ;
        RECT  28.30 7.10 29.00 11.00 ;
        RECT  0.00 11.00 30.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.45 ;
        RECT  6.50 2.00 7.20 4.40 ;
        RECT  11.05 2.00 11.75 4.85 ;
        RECT  15.15 2.00 16.75 3.15 ;
        RECT  16.05 2.00 16.75 4.90 ;
        RECT  18.20 2.00 18.90 3.25 ;
        RECT  24.05 2.00 24.75 3.95 ;
        RECT  28.30 2.00 29.00 4.45 ;
        RECT  0.00 0.00 30.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.15 3.95 5.20 4.45 ;
        RECT  7.85 9.60 9.70 9.95 ;
        RECT  0.45 3.75 0.95 9.90 ;
        RECT  0.45 3.75 1.15 4.45 ;
        RECT  0.45 8.10 1.15 9.90 ;
        RECT  3.50 6.85 4.20 7.55 ;
        RECT  0.45 7.05 4.20 7.55 ;
        RECT  4.70 3.75 4.85 9.90 ;
        RECT  4.15 8.15 4.85 9.90 ;
        RECT  4.70 3.75 5.05 8.65 ;
        RECT  4.15 3.75 5.05 4.45 ;
        RECT  4.70 3.95 5.20 8.65 ;
        RECT  4.15 8.15 5.20 8.65 ;
        RECT  8.15 8.10 8.55 10.30 ;
        RECT  7.85 8.10 8.55 9.95 ;
        RECT  7.85 3.75 9.20 4.50 ;
        RECT  8.70 3.75 9.20 6.35 ;
        RECT  8.70 5.65 9.55 6.35 ;
        RECT  8.15 9.60 9.70 10.30 ;
        RECT  9.70 4.20 10.55 4.90 ;
        RECT  9.70 8.00 10.40 9.00 ;
        RECT  10.05 4.20 10.55 6.05 ;
        RECT  11.50 6.65 12.20 7.35 ;
        RECT  4.70 6.85 12.20 7.35 ;
        RECT  10.05 5.55 13.35 6.05 ;
        RECT  12.35 3.20 12.85 6.05 ;
        RECT  12.85 5.55 13.35 8.50 ;
        RECT  9.70 8.00 13.35 8.50 ;
        RECT  12.85 6.70 13.55 7.40 ;
        RECT  13.40 4.20 14.10 4.90 ;
        RECT  13.40 4.40 14.55 4.90 ;
        RECT  14.05 4.20 14.10 9.70 ;
        RECT  13.40 9.00 14.10 9.70 ;
        RECT  13.85 3.00 14.55 3.70 ;
        RECT  12.35 3.20 14.55 3.70 ;
        RECT  14.05 4.40 14.55 9.50 ;
        RECT  13.40 9.00 14.55 9.50 ;
        RECT  15.30 5.45 16.00 6.15 ;
        RECT  14.05 6.70 16.95 7.20 ;
        RECT  16.25 6.70 16.95 7.40 ;
        RECT  15.30 5.45 17.95 5.95 ;
        RECT  17.45 4.35 17.95 9.70 ;
        RECT  17.45 9.00 18.25 9.70 ;
        RECT  18.55 4.15 19.25 4.85 ;
        RECT  17.45 4.35 19.25 4.85 ;
        RECT  20.70 3.30 21.40 4.00 ;
        RECT  20.70 3.45 22.60 4.00 ;
        RECT  21.55 7.20 22.10 10.50 ;
        RECT  21.40 8.75 22.10 10.50 ;
        RECT  22.10 3.45 22.60 7.90 ;
        RECT  21.55 7.20 22.60 7.90 ;
        RECT  23.60 4.45 24.30 5.15 ;
        RECT  24.40 5.70 25.10 6.40 ;
        RECT  22.10 5.90 25.10 6.40 ;
        RECT  25.40 3.25 26.10 3.95 ;
        RECT  23.60 4.45 26.10 4.95 ;
        RECT  25.60 3.25 26.10 10.50 ;
        RECT  25.40 7.40 26.10 10.50 ;
    END
END SDFRRX2
MACRO SDFRRX4
    CLASS CORE ;
    FOREIGN SDFRRX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 33.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  1.45 5.60 2.55 6.30 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END SD
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  18.45 7.05 19.15 8.40 ;
        RECT  19.85 6.70 20.75 7.60 ;
        RECT  20.25 5.45 20.75 7.60 ;
        RECT  18.45 7.05 20.75 7.60 ;
        RECT  20.90 5.25 21.60 5.95 ;
        RECT  20.25 5.45 21.60 5.95 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  31.10 2.50 31.80 4.10 ;
        RECT  31.30 2.50 31.80 10.50 ;
        RECT  31.10 5.35 31.80 10.50 ;
        RECT  30.95 5.35 31.95 6.35 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  28.40 2.50 28.90 10.50 ;
        RECT  28.40 2.50 29.10 4.10 ;
        RECT  28.40 8.10 29.10 10.50 ;
        RECT  28.25 5.35 29.15 6.35 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  6.50 8.10 7.20 11.00 ;
        RECT  11.05 9.00 11.75 11.00 ;
        RECT  15.75 7.90 16.45 11.00 ;
        RECT  19.05 8.90 19.75 11.00 ;
        RECT  24.05 7.40 24.75 11.00 ;
        RECT  27.05 8.10 27.75 11.00 ;
        RECT  29.75 8.10 30.45 11.00 ;
        RECT  32.45 8.10 33.15 11.00 ;
        RECT  0.00 11.00 33.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.45 ;
        RECT  6.50 2.00 7.20 4.40 ;
        RECT  11.05 2.00 11.75 4.85 ;
        RECT  15.15 2.00 16.75 3.15 ;
        RECT  16.05 2.00 16.75 4.90 ;
        RECT  18.20 2.00 18.90 3.25 ;
        RECT  24.05 2.00 24.75 3.95 ;
        RECT  27.05 2.00 27.75 4.10 ;
        RECT  29.75 2.00 30.45 4.10 ;
        RECT  32.45 2.00 33.15 4.10 ;
        RECT  0.00 0.00 33.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.15 3.95 5.20 4.45 ;
        RECT  7.85 9.60 9.70 9.95 ;
        RECT  0.45 3.75 0.95 9.90 ;
        RECT  0.45 3.75 1.15 4.45 ;
        RECT  0.45 8.10 1.15 9.90 ;
        RECT  3.50 6.85 4.20 7.55 ;
        RECT  0.45 7.05 4.20 7.55 ;
        RECT  4.70 3.75 4.85 9.90 ;
        RECT  4.15 8.15 4.85 9.90 ;
        RECT  4.70 3.75 5.05 8.65 ;
        RECT  4.15 3.75 5.05 4.45 ;
        RECT  4.70 3.95 5.20 8.65 ;
        RECT  4.15 8.15 5.20 8.65 ;
        RECT  8.15 8.10 8.55 10.30 ;
        RECT  7.85 8.10 8.55 9.95 ;
        RECT  7.85 3.75 9.20 4.50 ;
        RECT  8.70 3.75 9.20 6.35 ;
        RECT  8.70 5.65 9.55 6.35 ;
        RECT  8.15 9.60 9.70 10.30 ;
        RECT  9.70 4.20 10.55 4.90 ;
        RECT  9.70 8.00 10.40 9.00 ;
        RECT  10.05 4.20 10.55 6.05 ;
        RECT  11.50 6.65 12.20 7.35 ;
        RECT  4.70 6.85 12.20 7.35 ;
        RECT  10.05 5.55 13.35 6.05 ;
        RECT  12.35 3.20 12.85 6.05 ;
        RECT  12.85 5.55 13.35 8.50 ;
        RECT  9.70 8.00 13.35 8.50 ;
        RECT  12.85 6.70 13.55 7.40 ;
        RECT  13.40 4.20 14.10 4.90 ;
        RECT  13.40 4.40 14.55 4.90 ;
        RECT  14.05 4.20 14.10 9.70 ;
        RECT  13.40 9.00 14.10 9.70 ;
        RECT  13.85 3.00 14.55 3.70 ;
        RECT  12.35 3.20 14.55 3.70 ;
        RECT  14.05 4.40 14.55 9.50 ;
        RECT  13.40 9.00 14.55 9.50 ;
        RECT  15.30 5.45 16.00 6.15 ;
        RECT  14.05 6.70 16.95 7.20 ;
        RECT  16.25 6.70 16.95 7.40 ;
        RECT  15.30 5.45 17.95 5.95 ;
        RECT  17.45 4.35 17.95 9.70 ;
        RECT  17.45 9.00 18.25 9.70 ;
        RECT  18.55 4.15 19.25 4.85 ;
        RECT  17.45 4.35 19.25 4.85 ;
        RECT  20.70 3.30 21.40 4.00 ;
        RECT  20.70 3.45 22.60 4.00 ;
        RECT  21.55 7.20 22.10 10.50 ;
        RECT  21.40 8.75 22.10 10.50 ;
        RECT  22.10 3.45 22.60 7.90 ;
        RECT  21.55 7.20 22.60 7.90 ;
        RECT  23.60 4.45 24.30 5.15 ;
        RECT  24.40 5.70 25.10 6.40 ;
        RECT  22.10 5.90 25.10 6.40 ;
        RECT  25.40 3.25 26.10 3.95 ;
        RECT  23.60 4.45 26.70 4.95 ;
        RECT  25.60 3.25 26.10 10.10 ;
        RECT  25.40 7.40 26.10 10.10 ;
        RECT  25.60 4.45 26.70 5.15 ;
    END
END SDFRRX4
MACRO SDFRSX1
    CLASS CORE ;
    FOREIGN SDFRSX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 32.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  16.50 2.55 23.55 3.25 ;
        RECT  22.65 2.55 23.55 3.75 ;
        RECT  16.50 2.55 26.70 3.05 ;
        RECT  26.00 2.55 26.70 3.25 ;
        END
    END SN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  1.45 5.60 2.55 6.30 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END SD
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  28.35 2.65 29.05 4.30 ;
        RECT  28.35 7.25 29.05 9.75 ;
        RECT  28.35 3.80 30.15 4.30 ;
        RECT  29.65 3.80 30.15 7.75 ;
        RECT  28.35 7.25 30.15 7.75 ;
        RECT  29.65 5.35 30.55 6.35 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  31.05 2.65 31.75 3.35 ;
        RECT  31.25 2.65 31.75 9.75 ;
        RECT  31.05 7.95 31.75 9.75 ;
        RECT  30.95 7.95 31.95 8.95 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  6.50 8.10 7.20 11.00 ;
        RECT  11.05 8.85 11.75 11.00 ;
        RECT  16.80 8.20 17.50 11.00 ;
        RECT  19.30 9.55 20.00 11.00 ;
        RECT  24.15 9.30 24.85 11.00 ;
        RECT  26.85 9.30 27.55 11.00 ;
        RECT  29.70 8.25 30.40 11.00 ;
        RECT  0.00 11.00 32.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.45 ;
        RECT  6.50 2.00 7.20 4.40 ;
        RECT  11.05 2.00 11.75 4.85 ;
        RECT  15.50 2.00 16.00 4.25 ;
        RECT  16.90 3.75 17.60 4.95 ;
        RECT  15.50 3.75 20.60 4.25 ;
        RECT  19.90 3.75 20.60 5.45 ;
        RECT  25.55 3.75 26.25 5.45 ;
        RECT  24.60 4.70 26.25 5.45 ;
        RECT  27.35 2.00 27.85 4.25 ;
        RECT  25.55 3.75 27.85 4.25 ;
        RECT  29.70 2.00 30.40 3.30 ;
        RECT  0.00 0.00 32.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.15 3.95 5.20 4.45 ;
        RECT  23.95 6.05 29.15 6.50 ;
        RECT  7.85 9.60 9.70 9.95 ;
        RECT  0.45 3.75 0.95 9.90 ;
        RECT  0.45 3.75 1.15 4.45 ;
        RECT  0.45 8.10 1.15 9.90 ;
        RECT  3.50 6.85 4.20 7.55 ;
        RECT  0.45 7.05 4.20 7.55 ;
        RECT  4.70 3.75 4.85 9.90 ;
        RECT  4.15 8.15 4.85 9.90 ;
        RECT  4.70 3.75 5.05 8.65 ;
        RECT  4.15 3.75 5.05 4.45 ;
        RECT  4.70 3.95 5.20 8.65 ;
        RECT  4.15 8.15 5.20 8.65 ;
        RECT  8.15 8.10 8.55 10.30 ;
        RECT  7.85 8.10 8.55 9.95 ;
        RECT  7.85 3.75 9.20 4.50 ;
        RECT  8.70 3.75 9.20 6.35 ;
        RECT  8.70 5.65 9.55 6.35 ;
        RECT  8.15 9.60 9.70 10.30 ;
        RECT  9.70 4.20 10.55 4.90 ;
        RECT  9.70 7.85 10.40 8.90 ;
        RECT  10.05 4.20 10.55 6.05 ;
        RECT  11.50 6.65 12.20 7.35 ;
        RECT  4.70 6.85 12.20 7.35 ;
        RECT  10.05 5.55 13.20 6.05 ;
        RECT  12.70 3.20 12.85 8.35 ;
        RECT  12.35 3.20 12.85 6.05 ;
        RECT  12.70 5.55 13.20 8.35 ;
        RECT  9.70 7.85 13.20 8.35 ;
        RECT  12.70 6.70 13.55 7.40 ;
        RECT  13.40 4.20 14.55 4.90 ;
        RECT  13.85 3.00 14.55 3.70 ;
        RECT  12.35 3.20 14.55 3.70 ;
        RECT  14.05 4.20 14.55 9.50 ;
        RECT  13.40 8.80 15.00 9.50 ;
        RECT  16.35 5.65 17.05 6.35 ;
        RECT  17.35 6.90 18.05 7.60 ;
        RECT  14.05 7.10 18.05 7.60 ;
        RECT  18.40 4.75 19.10 6.15 ;
        RECT  16.35 5.65 19.10 6.15 ;
        RECT  18.60 4.75 19.10 8.85 ;
        RECT  18.15 8.10 19.10 8.85 ;
        RECT  22.25 4.75 22.50 10.05 ;
        RECT  21.80 7.30 22.50 10.05 ;
        RECT  22.25 4.75 22.75 7.80 ;
        RECT  22.25 4.75 22.95 5.45 ;
        RECT  23.95 6.00 24.65 6.70 ;
        RECT  25.50 8.30 26.20 9.95 ;
        RECT  26.15 7.10 26.85 7.80 ;
        RECT  21.80 7.30 26.85 7.80 ;
        RECT  27.35 6.00 27.85 8.80 ;
        RECT  25.50 8.30 27.85 8.80 ;
        RECT  27.90 4.80 28.60 6.75 ;
        RECT  23.95 6.00 28.60 6.50 ;
        RECT  27.35 6.05 29.15 6.75 ;
    END
END SDFRSX1
MACRO SDFRSX2
    CLASS CORE ;
    FOREIGN SDFRSX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 32.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  16.50 2.55 23.55 3.25 ;
        RECT  22.65 2.55 23.55 3.75 ;
        RECT  16.50 2.55 26.70 3.05 ;
        RECT  26.00 2.55 26.70 3.25 ;
        END
    END SN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  1.45 5.60 2.55 6.30 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END SD
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  28.35 2.65 29.05 4.30 ;
        RECT  28.35 7.25 29.05 10.50 ;
        RECT  28.35 3.80 30.15 4.30 ;
        RECT  29.65 3.80 30.15 7.75 ;
        RECT  28.35 7.25 30.15 7.75 ;
        RECT  29.65 5.35 30.55 6.35 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  31.05 2.65 31.75 3.35 ;
        RECT  31.25 2.65 31.75 10.50 ;
        RECT  31.05 7.95 31.75 10.50 ;
        RECT  30.95 7.95 31.95 8.95 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  6.50 8.10 7.20 11.00 ;
        RECT  11.05 8.85 11.75 11.00 ;
        RECT  16.80 8.20 17.50 11.00 ;
        RECT  19.30 9.55 20.00 11.00 ;
        RECT  24.15 9.30 24.85 11.00 ;
        RECT  26.85 9.30 27.55 11.00 ;
        RECT  29.70 8.25 30.40 11.00 ;
        RECT  0.00 11.00 32.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.45 ;
        RECT  6.50 2.00 7.20 4.40 ;
        RECT  11.05 2.00 11.75 4.85 ;
        RECT  15.50 2.00 16.00 4.25 ;
        RECT  16.90 3.75 17.60 4.95 ;
        RECT  15.50 3.75 20.60 4.25 ;
        RECT  19.90 3.75 20.60 5.45 ;
        RECT  25.55 3.75 26.25 5.45 ;
        RECT  24.60 4.70 26.25 5.45 ;
        RECT  27.35 2.00 27.85 4.25 ;
        RECT  25.55 3.75 27.85 4.25 ;
        RECT  29.70 2.00 30.40 3.30 ;
        RECT  0.00 0.00 32.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.15 3.95 5.20 4.45 ;
        RECT  23.95 6.05 29.15 6.50 ;
        RECT  7.85 9.60 9.70 9.95 ;
        RECT  0.45 3.75 0.95 9.90 ;
        RECT  0.45 3.75 1.15 4.45 ;
        RECT  0.45 8.10 1.15 9.90 ;
        RECT  3.50 6.85 4.20 7.55 ;
        RECT  0.45 7.05 4.20 7.55 ;
        RECT  4.70 3.75 4.85 9.90 ;
        RECT  4.15 8.15 4.85 9.90 ;
        RECT  4.70 3.75 5.05 8.65 ;
        RECT  4.15 3.75 5.05 4.45 ;
        RECT  4.70 3.95 5.20 8.65 ;
        RECT  4.15 8.15 5.20 8.65 ;
        RECT  8.15 8.10 8.55 10.30 ;
        RECT  7.85 8.10 8.55 9.95 ;
        RECT  7.85 3.75 9.20 4.50 ;
        RECT  8.70 3.75 9.20 6.35 ;
        RECT  8.70 5.65 9.55 6.35 ;
        RECT  8.15 9.60 9.70 10.30 ;
        RECT  9.70 4.20 10.55 4.90 ;
        RECT  9.70 7.85 10.40 8.90 ;
        RECT  10.05 4.20 10.55 6.05 ;
        RECT  11.50 6.65 12.20 7.35 ;
        RECT  4.70 6.85 12.20 7.35 ;
        RECT  10.05 5.55 13.20 6.05 ;
        RECT  12.70 3.20 12.85 8.35 ;
        RECT  12.35 3.20 12.85 6.05 ;
        RECT  12.70 5.55 13.20 8.35 ;
        RECT  9.70 7.85 13.20 8.35 ;
        RECT  12.70 6.70 13.55 7.40 ;
        RECT  13.40 4.20 14.55 4.90 ;
        RECT  13.85 3.00 14.55 3.70 ;
        RECT  12.35 3.20 14.55 3.70 ;
        RECT  14.05 4.20 14.55 9.50 ;
        RECT  13.40 8.80 15.00 9.50 ;
        RECT  16.35 5.65 17.05 6.35 ;
        RECT  17.35 6.90 18.05 7.60 ;
        RECT  14.05 7.10 18.05 7.60 ;
        RECT  18.40 4.75 19.10 6.15 ;
        RECT  16.35 5.65 19.10 6.15 ;
        RECT  18.60 4.75 19.10 8.85 ;
        RECT  18.15 8.10 19.10 8.85 ;
        RECT  22.25 4.75 22.50 10.05 ;
        RECT  21.80 7.30 22.50 10.05 ;
        RECT  22.25 4.75 22.75 7.80 ;
        RECT  22.25 4.75 22.95 5.45 ;
        RECT  23.95 6.00 24.65 6.70 ;
        RECT  25.50 8.30 26.20 9.95 ;
        RECT  26.15 7.10 26.85 7.80 ;
        RECT  21.80 7.30 26.85 7.80 ;
        RECT  27.35 6.00 27.85 8.80 ;
        RECT  25.50 8.30 27.85 8.80 ;
        RECT  27.90 4.80 28.60 6.75 ;
        RECT  23.95 6.00 28.60 6.50 ;
        RECT  27.35 6.05 29.15 6.75 ;
    END
END SDFRSX2
MACRO SDFRSX4
    CLASS CORE ;
    FOREIGN SDFRSX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 35.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  16.50 2.55 23.55 3.25 ;
        RECT  22.65 2.55 23.55 3.75 ;
        RECT  16.50 2.55 26.70 3.05 ;
        RECT  26.00 2.55 26.70 3.25 ;
        END
    END SN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  1.45 5.60 2.55 6.30 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END SD
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  29.80 2.50 30.30 10.50 ;
        RECT  29.80 2.50 30.50 4.10 ;
        RECT  29.80 8.10 30.50 10.50 ;
        RECT  29.65 5.35 30.55 6.35 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  32.50 2.50 33.20 4.10 ;
        RECT  32.70 2.50 33.20 10.50 ;
        RECT  32.50 5.35 33.20 10.50 ;
        RECT  32.35 5.35 33.35 6.35 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  6.50 8.10 7.20 11.00 ;
        RECT  11.05 8.85 11.75 11.00 ;
        RECT  16.80 8.20 17.50 11.00 ;
        RECT  19.30 9.55 20.00 11.00 ;
        RECT  24.15 9.30 24.85 11.00 ;
        RECT  26.85 9.30 27.55 11.00 ;
        RECT  28.45 8.10 29.15 11.00 ;
        RECT  31.15 8.10 31.85 11.00 ;
        RECT  33.85 8.10 34.55 11.00 ;
        RECT  0.00 11.00 35.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.45 ;
        RECT  6.50 2.00 7.20 4.40 ;
        RECT  11.05 2.00 11.75 4.85 ;
        RECT  15.50 2.00 16.00 4.25 ;
        RECT  16.90 3.75 17.60 4.95 ;
        RECT  15.50 3.75 20.60 4.25 ;
        RECT  19.90 3.75 20.60 5.45 ;
        RECT  25.55 3.75 26.25 5.45 ;
        RECT  24.60 4.70 26.25 5.45 ;
        RECT  28.30 2.00 29.00 4.25 ;
        RECT  25.55 3.75 29.00 4.25 ;
        RECT  31.15 2.00 31.85 4.10 ;
        RECT  33.85 2.00 34.55 4.10 ;
        RECT  0.00 0.00 35.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.15 3.95 5.20 4.45 ;
        RECT  7.85 9.60 9.70 9.95 ;
        RECT  0.45 3.75 0.95 9.90 ;
        RECT  0.45 3.75 1.15 4.45 ;
        RECT  0.45 8.10 1.15 9.90 ;
        RECT  3.50 6.85 4.20 7.55 ;
        RECT  0.45 7.05 4.20 7.55 ;
        RECT  4.70 3.75 4.85 9.90 ;
        RECT  4.15 8.15 4.85 9.90 ;
        RECT  4.70 3.75 5.05 8.65 ;
        RECT  4.15 3.75 5.05 4.45 ;
        RECT  4.70 3.95 5.20 8.65 ;
        RECT  4.15 8.15 5.20 8.65 ;
        RECT  8.15 8.10 8.55 10.30 ;
        RECT  7.85 8.10 8.55 9.95 ;
        RECT  7.85 3.75 9.20 4.50 ;
        RECT  8.70 3.75 9.20 6.35 ;
        RECT  8.70 5.65 9.55 6.35 ;
        RECT  8.15 9.60 9.70 10.30 ;
        RECT  9.70 4.20 10.55 4.90 ;
        RECT  9.70 7.85 10.40 8.90 ;
        RECT  10.05 4.20 10.55 6.05 ;
        RECT  11.50 6.65 12.20 7.35 ;
        RECT  4.70 6.85 12.20 7.35 ;
        RECT  10.05 5.55 13.20 6.05 ;
        RECT  12.70 3.20 12.85 8.35 ;
        RECT  12.35 3.20 12.85 6.05 ;
        RECT  12.70 5.55 13.20 8.35 ;
        RECT  9.70 7.85 13.20 8.35 ;
        RECT  12.70 6.70 13.55 7.40 ;
        RECT  13.40 4.20 14.55 4.90 ;
        RECT  13.85 3.00 14.55 3.70 ;
        RECT  12.35 3.20 14.55 3.70 ;
        RECT  14.05 4.20 14.55 9.50 ;
        RECT  13.40 8.80 15.00 9.50 ;
        RECT  16.35 5.65 17.05 6.35 ;
        RECT  17.35 6.90 18.05 7.60 ;
        RECT  14.05 7.10 18.05 7.60 ;
        RECT  18.40 4.75 19.10 6.15 ;
        RECT  16.35 5.65 19.10 6.15 ;
        RECT  18.60 4.75 19.10 8.85 ;
        RECT  18.15 8.10 19.10 8.85 ;
        RECT  22.25 4.75 22.50 10.05 ;
        RECT  21.80 7.30 22.50 10.05 ;
        RECT  22.25 4.75 22.75 7.80 ;
        RECT  22.25 4.75 22.95 5.45 ;
        RECT  23.95 6.00 24.65 6.70 ;
        RECT  25.50 8.30 26.20 9.95 ;
        RECT  26.15 7.10 26.85 7.80 ;
        RECT  21.80 7.30 26.85 7.80 ;
        RECT  27.35 6.00 27.85 8.80 ;
        RECT  25.50 8.30 27.85 8.80 ;
        RECT  23.95 6.00 29.15 6.50 ;
        RECT  28.45 4.80 28.60 6.70 ;
        RECT  27.90 4.80 28.60 6.50 ;
        RECT  28.45 6.00 29.15 6.70 ;
    END
END SDFRSX4
MACRO SDFRX1
    CLASS CORE ;
    FOREIGN SDFRX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 28.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  1.45 5.60 2.55 6.30 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END SD
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  26.85 3.75 27.55 4.45 ;
        RECT  27.05 3.75 27.55 8.85 ;
        RECT  26.85 7.15 27.55 8.85 ;
        RECT  26.85 5.40 27.75 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  24.15 3.75 24.85 4.45 ;
        RECT  24.30 3.75 24.85 8.85 ;
        RECT  24.15 7.15 24.85 8.85 ;
        RECT  24.05 5.40 24.95 6.30 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  21.45 8.60 22.30 9.10 ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  6.50 8.10 7.20 11.00 ;
        RECT  11.05 8.85 11.75 11.00 ;
        RECT  15.75 7.90 16.45 11.00 ;
        RECT  15.00 10.45 16.60 11.00 ;
        RECT  17.95 10.40 18.65 11.00 ;
        RECT  21.25 7.40 21.95 8.15 ;
        RECT  21.80 7.40 21.95 11.00 ;
        RECT  21.45 7.40 21.95 9.10 ;
        RECT  21.80 8.60 22.30 11.00 ;
        RECT  21.80 10.15 23.50 11.00 ;
        RECT  25.50 7.15 26.20 11.00 ;
        RECT  24.30 10.70 27.55 11.00 ;
        RECT  0.00 11.00 28.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.45 ;
        RECT  6.50 2.00 7.20 4.40 ;
        RECT  11.05 2.00 11.75 4.85 ;
        RECT  15.80 2.00 16.55 4.90 ;
        RECT  21.25 2.00 21.95 3.95 ;
        RECT  25.50 2.00 26.20 4.45 ;
        RECT  0.00 0.00 28.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.15 3.95 5.20 4.45 ;
        RECT  7.85 9.60 9.70 9.95 ;
        RECT  0.45 3.75 0.95 9.90 ;
        RECT  0.45 3.75 1.15 4.45 ;
        RECT  0.45 8.10 1.15 9.90 ;
        RECT  3.50 6.85 4.20 7.55 ;
        RECT  0.45 7.05 4.20 7.55 ;
        RECT  4.70 3.75 4.85 9.90 ;
        RECT  4.15 8.15 4.85 9.90 ;
        RECT  4.70 3.75 5.05 8.65 ;
        RECT  4.15 3.75 5.05 4.45 ;
        RECT  4.70 3.95 5.20 8.65 ;
        RECT  4.15 8.15 5.20 8.65 ;
        RECT  8.15 8.10 8.55 10.30 ;
        RECT  7.85 8.10 8.55 9.95 ;
        RECT  7.85 3.75 9.20 4.50 ;
        RECT  8.70 3.75 9.20 6.35 ;
        RECT  8.70 5.65 9.55 6.35 ;
        RECT  8.15 9.60 9.70 10.30 ;
        RECT  9.70 4.20 10.55 4.90 ;
        RECT  9.70 7.85 10.40 8.90 ;
        RECT  10.05 4.20 10.55 6.05 ;
        RECT  11.50 6.65 12.20 7.35 ;
        RECT  4.70 6.85 12.20 7.35 ;
        RECT  10.05 5.55 13.20 6.05 ;
        RECT  12.70 3.20 12.85 8.35 ;
        RECT  12.35 3.20 12.85 6.05 ;
        RECT  12.70 5.55 13.20 8.35 ;
        RECT  9.70 7.85 13.20 8.35 ;
        RECT  12.70 6.70 13.55 7.40 ;
        RECT  13.40 4.20 14.10 4.90 ;
        RECT  13.40 4.40 14.55 4.90 ;
        RECT  14.05 4.20 14.10 9.50 ;
        RECT  13.40 8.80 14.10 9.50 ;
        RECT  13.85 3.00 14.55 3.70 ;
        RECT  12.35 3.20 14.55 3.70 ;
        RECT  14.05 4.40 14.55 9.30 ;
        RECT  13.40 8.80 14.55 9.30 ;
        RECT  15.30 5.45 16.00 6.15 ;
        RECT  14.05 6.70 16.95 7.20 ;
        RECT  16.25 6.70 16.95 7.40 ;
        RECT  17.25 4.15 17.95 4.85 ;
        RECT  15.30 5.45 17.95 5.95 ;
        RECT  17.45 4.15 17.95 8.60 ;
        RECT  17.25 7.90 17.95 8.60 ;
        RECT  18.90 3.30 19.60 4.00 ;
        RECT  19.10 3.30 19.60 10.15 ;
        RECT  19.10 9.65 21.00 10.15 ;
        RECT  20.30 9.65 21.00 10.35 ;
        RECT  20.80 4.45 21.50 5.15 ;
        RECT  21.60 5.70 22.30 6.40 ;
        RECT  19.10 5.90 22.30 6.40 ;
        RECT  22.60 3.25 23.30 3.95 ;
        RECT  20.80 4.45 23.30 4.95 ;
        RECT  22.60 7.40 23.30 8.15 ;
        RECT  22.80 3.25 23.30 9.65 ;
        RECT  22.80 8.95 23.65 9.65 ;
    END
END SDFRX1
MACRO SDFRX2
    CLASS CORE ;
    FOREIGN SDFRX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 28.00 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  1.45 5.60 2.55 6.30 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END SD
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  26.85 2.75 27.55 4.45 ;
        RECT  27.05 2.75 27.55 10.50 ;
        RECT  26.85 7.10 27.55 10.50 ;
        RECT  26.85 5.40 27.75 6.30 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  24.15 2.75 24.85 4.45 ;
        RECT  24.30 2.75 24.85 9.60 ;
        RECT  24.15 7.10 24.85 9.60 ;
        RECT  24.05 5.40 24.95 6.30 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  21.45 8.60 22.30 9.10 ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  6.50 8.10 7.20 11.00 ;
        RECT  11.05 8.85 11.75 11.00 ;
        RECT  15.75 7.90 16.45 11.00 ;
        RECT  15.00 10.45 16.60 11.00 ;
        RECT  17.95 10.40 18.65 11.00 ;
        RECT  21.25 7.40 21.95 8.15 ;
        RECT  21.80 7.40 21.95 11.00 ;
        RECT  21.45 7.40 21.95 9.10 ;
        RECT  21.80 8.60 22.30 11.00 ;
        RECT  21.80 10.20 23.50 11.00 ;
        RECT  17.95 10.85 23.50 11.00 ;
        RECT  25.50 7.10 26.20 11.00 ;
        RECT  0.00 11.00 28.00 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.45 ;
        RECT  6.50 2.00 7.20 4.40 ;
        RECT  11.05 2.00 11.75 4.85 ;
        RECT  15.80 2.00 16.55 4.90 ;
        RECT  21.25 2.00 21.95 3.95 ;
        RECT  25.50 2.00 26.20 4.45 ;
        RECT  0.00 0.00 28.00 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.15 3.95 5.20 4.45 ;
        RECT  7.85 9.60 9.70 9.95 ;
        RECT  0.45 3.75 0.95 9.90 ;
        RECT  0.45 3.75 1.15 4.45 ;
        RECT  0.45 8.10 1.15 9.90 ;
        RECT  3.50 6.85 4.20 7.55 ;
        RECT  0.45 7.05 4.20 7.55 ;
        RECT  4.70 3.75 4.85 9.90 ;
        RECT  4.15 8.15 4.85 9.90 ;
        RECT  4.70 3.75 5.05 8.65 ;
        RECT  4.15 3.75 5.05 4.45 ;
        RECT  4.70 3.95 5.20 8.65 ;
        RECT  4.15 8.15 5.20 8.65 ;
        RECT  8.15 8.10 8.55 10.30 ;
        RECT  7.85 8.10 8.55 9.95 ;
        RECT  7.85 3.75 9.20 4.50 ;
        RECT  8.70 3.75 9.20 6.35 ;
        RECT  8.70 5.65 9.55 6.35 ;
        RECT  8.15 9.60 9.70 10.30 ;
        RECT  9.70 4.20 10.55 4.90 ;
        RECT  9.70 7.85 10.40 8.90 ;
        RECT  10.05 4.20 10.55 6.05 ;
        RECT  11.50 6.65 12.20 7.35 ;
        RECT  4.70 6.85 12.20 7.35 ;
        RECT  10.05 5.55 13.20 6.05 ;
        RECT  12.70 3.20 12.85 8.35 ;
        RECT  12.35 3.20 12.85 6.05 ;
        RECT  12.70 5.55 13.20 8.35 ;
        RECT  9.70 7.85 13.20 8.35 ;
        RECT  12.70 6.70 13.55 7.40 ;
        RECT  13.40 4.20 14.10 4.90 ;
        RECT  13.40 4.40 14.55 4.90 ;
        RECT  14.05 4.20 14.10 9.50 ;
        RECT  13.40 8.80 14.10 9.50 ;
        RECT  13.85 3.00 14.55 3.70 ;
        RECT  12.35 3.20 14.55 3.70 ;
        RECT  14.05 4.40 14.55 9.30 ;
        RECT  13.40 8.80 14.55 9.30 ;
        RECT  15.30 5.45 16.00 6.15 ;
        RECT  14.05 6.70 16.95 7.20 ;
        RECT  16.25 6.70 16.95 7.40 ;
        RECT  17.25 4.15 17.95 4.85 ;
        RECT  15.30 5.45 17.95 5.95 ;
        RECT  17.45 4.15 17.95 8.60 ;
        RECT  17.25 7.90 17.95 8.60 ;
        RECT  18.90 3.30 19.60 4.00 ;
        RECT  19.10 3.30 19.60 10.15 ;
        RECT  19.10 9.65 21.00 10.15 ;
        RECT  20.30 9.65 21.00 10.35 ;
        RECT  20.80 4.45 21.50 5.15 ;
        RECT  21.60 5.70 22.30 6.40 ;
        RECT  19.10 5.90 22.30 6.40 ;
        RECT  22.60 3.25 23.30 3.95 ;
        RECT  20.80 4.45 23.30 4.95 ;
        RECT  22.60 7.40 23.30 8.15 ;
        RECT  22.80 3.25 23.30 9.65 ;
        RECT  22.80 8.95 23.65 9.65 ;
    END
END SDFRX2
MACRO SDFRX4
    CLASS CORE ;
    FOREIGN SDFRX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 30.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.10 ;
        PORT
        LAYER M1M ;
        RECT  1.65 5.40 2.55 6.30 ;
        RECT  1.45 5.60 2.55 6.30 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  3.05 5.40 3.95 6.30 ;
        END
    END SD
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  28.30 2.90 29.00 4.50 ;
        RECT  28.50 2.90 29.00 10.50 ;
        RECT  28.30 5.35 29.00 10.50 ;
        RECT  28.15 5.35 29.15 6.35 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  25.60 2.90 26.10 10.50 ;
        RECT  25.60 2.90 26.30 4.50 ;
        RECT  25.60 7.10 26.30 10.50 ;
        RECT  25.45 5.35 26.35 6.35 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  5.85 5.40 6.75 6.30 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  7.25 5.40 8.15 6.30 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 8.10 2.50 11.00 ;
        RECT  6.50 8.10 7.20 11.00 ;
        RECT  11.05 8.85 11.75 11.00 ;
        RECT  15.75 7.90 16.45 11.00 ;
        RECT  15.00 10.45 16.60 11.00 ;
        RECT  17.90 10.40 18.60 11.00 ;
        RECT  21.25 7.40 21.95 8.15 ;
        RECT  21.45 7.40 21.95 11.00 ;
        RECT  21.45 10.15 23.45 11.00 ;
        RECT  24.25 7.10 24.95 11.00 ;
        RECT  26.95 7.10 27.65 11.00 ;
        RECT  29.65 7.10 30.35 11.00 ;
        RECT  0.00 11.00 30.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 2.00 2.50 4.45 ;
        RECT  6.50 2.00 7.20 4.40 ;
        RECT  11.05 2.00 11.75 4.85 ;
        RECT  15.80 2.00 16.55 4.90 ;
        RECT  21.25 2.00 21.95 3.95 ;
        RECT  24.25 2.00 24.95 4.50 ;
        RECT  26.95 2.00 27.65 4.50 ;
        RECT  29.65 2.00 30.35 4.50 ;
        RECT  0.00 0.00 30.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  4.15 3.95 5.20 4.45 ;
        RECT  7.85 9.60 9.70 9.95 ;
        RECT  0.45 3.75 0.95 9.90 ;
        RECT  0.45 3.75 1.15 4.45 ;
        RECT  0.45 8.10 1.15 9.90 ;
        RECT  3.50 6.85 4.20 7.55 ;
        RECT  0.45 7.05 4.20 7.55 ;
        RECT  4.70 3.75 4.85 9.90 ;
        RECT  4.15 8.15 4.85 9.90 ;
        RECT  4.70 3.75 5.05 8.65 ;
        RECT  4.15 3.75 5.05 4.45 ;
        RECT  4.70 3.95 5.20 8.65 ;
        RECT  4.15 8.15 5.20 8.65 ;
        RECT  8.15 8.10 8.55 10.30 ;
        RECT  7.85 8.10 8.55 9.95 ;
        RECT  7.85 3.75 9.20 4.50 ;
        RECT  8.70 3.75 9.20 6.35 ;
        RECT  8.70 5.65 9.55 6.35 ;
        RECT  8.15 9.60 9.70 10.30 ;
        RECT  9.70 4.20 10.55 4.90 ;
        RECT  9.70 7.85 10.40 8.90 ;
        RECT  10.05 4.20 10.55 6.05 ;
        RECT  11.50 6.65 12.20 7.35 ;
        RECT  4.70 6.85 12.20 7.35 ;
        RECT  10.05 5.55 13.20 6.05 ;
        RECT  12.70 3.20 12.85 8.35 ;
        RECT  12.35 3.20 12.85 6.05 ;
        RECT  12.70 5.55 13.20 8.35 ;
        RECT  9.70 7.85 13.20 8.35 ;
        RECT  12.70 6.70 13.55 7.40 ;
        RECT  13.40 4.20 14.10 4.90 ;
        RECT  13.40 4.40 14.55 4.90 ;
        RECT  14.05 4.20 14.10 9.50 ;
        RECT  13.40 8.80 14.10 9.50 ;
        RECT  13.85 3.00 14.55 3.70 ;
        RECT  12.35 3.20 14.55 3.70 ;
        RECT  14.05 4.40 14.55 9.30 ;
        RECT  13.40 8.80 14.55 9.30 ;
        RECT  15.30 5.45 16.00 6.15 ;
        RECT  14.05 6.70 16.95 7.20 ;
        RECT  16.25 6.70 16.95 7.40 ;
        RECT  17.25 4.15 17.95 4.85 ;
        RECT  15.30 5.45 17.95 5.95 ;
        RECT  17.45 4.15 17.95 8.60 ;
        RECT  17.25 7.90 17.95 8.60 ;
        RECT  18.90 3.30 19.60 4.00 ;
        RECT  19.10 3.30 19.60 10.15 ;
        RECT  19.10 9.65 20.95 10.15 ;
        RECT  20.25 9.65 20.95 10.35 ;
        RECT  20.80 4.45 21.50 5.15 ;
        RECT  21.60 5.70 22.30 6.40 ;
        RECT  19.10 5.90 22.30 6.40 ;
        RECT  22.60 3.25 23.30 3.95 ;
        RECT  20.80 4.45 23.75 4.95 ;
        RECT  22.60 7.40 23.30 8.15 ;
        RECT  22.80 3.25 23.30 9.65 ;
        RECT  22.80 8.95 23.65 9.65 ;
        RECT  22.80 4.45 23.75 5.15 ;
    END
END SDFRX4
MACRO SIGNALHOLD
    CLASS CORE ;
    FOREIGN SIGNALHOLD 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SIG
        DIRECTION INOUT ;
        PORT
        LAYER M1M ;
        RECT  0.45 3.75 0.95 8.85 ;
        RECT  0.45 3.75 1.15 4.55 ;
        RECT  0.45 7.15 1.15 8.85 ;
        RECT  0.45 4.05 8.15 4.55 ;
        RECT  7.25 4.05 8.15 5.05 ;
        END
    END SIG
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.60 9.85 2.30 11.00 ;
        RECT  7.05 8.45 8.90 9.15 ;
        RECT  8.40 8.45 8.90 11.00 ;
        RECT  8.40 10.35 9.25 11.00 ;
        RECT  0.00 11.00 9.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  3.85 2.00 6.25 3.30 ;
        RECT  7.30 2.00 8.00 3.35 ;
        RECT  0.00 0.00 9.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  1.65 5.95 3.25 6.70 ;
        RECT  2.75 5.95 3.25 7.60 ;
        RECT  2.75 7.10 9.15 7.60 ;
        RECT  8.65 2.65 9.15 7.80 ;
        RECT  7.05 7.10 9.15 7.80 ;
        RECT  8.65 2.65 9.35 3.35 ;
    END
END SIGNALHOLD
MACRO SJKRRX1
    CLASS CORE ;
    FOREIGN SJKRRX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 44.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  28.25 5.40 29.15 6.30 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  26.85 5.40 27.75 6.30 ;
        END
    END SD
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  9.50 3.00 18.90 3.25 ;
        RECT  15.65 2.55 16.55 3.70 ;
        RECT  9.50 2.55 16.55 3.25 ;
        RECT  15.65 3.00 18.90 3.70 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M2M ;
        RECT  21.40 3.45 22.00 9.00 ;
        RECT  21.30 3.45 22.10 4.25 ;
        RECT  21.30 7.90 22.10 9.00 ;
        LAYER M1M ;
        RECT  21.35 3.10 22.05 4.30 ;
        RECT  21.35 8.00 22.05 9.75 ;
        RECT  21.25 3.40 22.15 4.30 ;
        RECT  21.25 8.00 22.15 8.90 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  24.05 3.10 24.75 3.80 ;
        RECT  24.25 3.10 24.75 9.75 ;
        RECT  24.05 7.95 24.75 9.75 ;
        RECT  24.05 7.95 24.95 8.95 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  40.85 5.40 41.75 6.30 ;
        RECT  40.30 5.60 41.75 6.30 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  42.25 5.40 43.15 6.30 ;
        END
    END J
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.25 6.65 2.55 7.35 ;
        RECT  1.65 6.65 2.55 7.65 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.30 2.50 11.00 ;
        RECT  4.05 7.95 4.75 11.00 ;
        RECT  9.80 8.10 10.50 11.00 ;
        RECT  12.30 9.55 13.00 11.00 ;
        RECT  17.15 9.05 17.85 11.00 ;
        RECT  19.85 9.15 20.55 11.00 ;
        RECT  22.70 8.25 23.40 11.00 ;
        RECT  27.20 7.10 27.90 11.00 ;
        RECT  39.40 7.80 40.10 11.00 ;
        RECT  42.25 7.10 42.95 11.00 ;
        RECT  0.00 11.00 44.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.90 2.00 1.70 3.20 ;
        RECT  4.05 2.00 4.75 4.85 ;
        RECT  8.50 2.00 9.00 4.25 ;
        RECT  9.90 3.75 10.60 4.95 ;
        RECT  8.50 3.75 13.60 4.25 ;
        RECT  12.90 3.75 13.60 5.40 ;
        RECT  17.60 4.65 19.25 5.40 ;
        RECT  19.40 2.00 19.90 5.15 ;
        RECT  17.60 4.65 19.90 5.15 ;
        RECT  22.70 2.00 23.40 3.75 ;
        RECT  27.20 2.00 27.90 4.45 ;
        RECT  34.20 2.00 34.90 4.15 ;
        RECT  42.25 2.00 42.95 4.45 ;
        RECT  0.00 0.00 44.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.25 5.35 0.75 10.25 ;
        RECT  0.25 9.55 1.15 10.25 ;
        RECT  1.00 3.80 1.80 5.85 ;
        RECT  0.25 5.35 1.80 5.85 ;
        RECT  2.70 4.20 3.55 4.90 ;
        RECT  3.05 4.20 3.55 8.85 ;
        RECT  2.70 8.15 3.55 8.85 ;
        RECT  3.05 5.55 6.35 6.05 ;
        RECT  5.35 3.20 5.85 6.05 ;
        RECT  5.85 5.55 6.35 7.40 ;
        RECT  5.85 6.70 6.55 7.40 ;
        RECT  6.40 4.20 7.55 4.90 ;
        RECT  6.85 3.00 7.55 3.70 ;
        RECT  5.35 3.20 7.55 3.70 ;
        RECT  7.05 4.20 7.55 9.25 ;
        RECT  6.40 8.55 8.00 9.25 ;
        RECT  9.35 5.65 10.05 6.35 ;
        RECT  10.35 6.90 11.05 7.60 ;
        RECT  7.05 7.10 11.05 7.60 ;
        RECT  11.40 4.75 12.10 6.15 ;
        RECT  9.35 5.65 12.10 6.15 ;
        RECT  11.60 4.75 12.10 8.85 ;
        RECT  11.15 8.10 12.10 8.85 ;
        RECT  15.25 4.70 15.50 9.85 ;
        RECT  14.80 7.15 15.50 9.85 ;
        RECT  15.25 4.70 15.75 7.65 ;
        RECT  15.25 4.70 15.95 5.40 ;
        RECT  16.95 5.95 17.65 6.70 ;
        RECT  18.50 8.15 19.20 9.85 ;
        RECT  19.00 6.95 19.70 7.65 ;
        RECT  14.80 7.15 19.70 7.65 ;
        RECT  16.95 5.95 20.70 6.45 ;
        RECT  20.20 5.75 20.70 8.65 ;
        RECT  18.50 8.15 20.70 8.65 ;
        RECT  20.90 4.75 21.60 6.25 ;
        RECT  20.20 5.75 23.75 6.25 ;
        RECT  23.05 5.55 23.75 6.25 ;
        RECT  16.95 5.95 23.75 6.25 ;
        RECT  25.50 2.55 26.35 3.25 ;
        RECT  25.80 2.55 26.35 8.90 ;
        RECT  25.80 3.75 26.55 4.45 ;
        RECT  25.80 7.10 26.60 8.90 ;
        RECT  28.55 3.75 29.25 4.45 ;
        RECT  28.55 7.10 29.25 8.90 ;
        RECT  28.55 3.95 30.15 4.45 ;
        RECT  29.65 3.95 30.15 7.60 ;
        RECT  28.55 7.10 30.15 7.60 ;
        RECT  30.20 9.75 30.90 10.45 ;
        RECT  30.65 4.60 31.35 5.30 ;
        RECT  31.50 6.80 32.00 9.45 ;
        RECT  31.30 7.75 32.00 9.45 ;
        RECT  31.65 3.70 32.35 5.10 ;
        RECT  32.65 7.80 33.35 10.45 ;
        RECT  30.20 9.95 33.35 10.45 ;
        RECT  34.00 6.80 34.70 10.45 ;
        RECT  35.35 7.80 36.05 10.45 ;
        RECT  31.50 6.80 37.20 7.30 ;
        RECT  36.70 6.80 37.20 9.45 ;
        RECT  36.70 7.75 37.40 9.45 ;
        RECT  37.40 5.60 38.10 6.30 ;
        RECT  29.65 5.80 38.10 6.30 ;
        RECT  37.70 3.45 38.20 5.10 ;
        RECT  30.65 4.60 38.20 5.10 ;
        RECT  38.05 7.80 38.75 10.45 ;
        RECT  38.25 6.80 38.75 10.45 ;
        RECT  35.35 9.95 38.75 10.45 ;
        RECT  37.70 3.45 39.30 4.15 ;
        RECT  38.25 6.80 41.25 7.30 ;
        RECT  40.75 6.80 41.25 10.50 ;
        RECT  40.75 7.80 41.45 10.50 ;
        RECT  43.65 3.75 44.15 10.50 ;
        RECT  43.65 3.75 44.35 4.45 ;
        RECT  43.65 7.10 44.35 10.50 ;
        RECT  43.65 9.80 44.50 10.50 ;
        LAYER V1M ;
        RECT  21.20 7.95 22.20 8.95 ;
        RECT  21.20 4.05 22.20 5.05 ;
        RECT  21.20 2.75 22.20 3.75 ;
    END
END SJKRRX1
MACRO SJKRRX2
    CLASS CORE ;
    FOREIGN SJKRRX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 44.80 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  28.25 5.40 29.15 6.30 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  26.85 5.40 27.75 6.30 ;
        END
    END SD
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  9.50 2.55 10.20 3.25 ;
        RECT  15.65 2.70 16.55 3.70 ;
        RECT  17.15 2.55 17.85 3.25 ;
        RECT  9.50 2.70 17.85 3.25 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M2M ;
        RECT  21.40 4.10 22.00 9.00 ;
        RECT  21.30 4.10 22.10 4.90 ;
        RECT  21.30 7.90 22.10 9.00 ;
        LAYER M1M ;
        RECT  21.35 2.75 22.05 4.95 ;
        RECT  21.35 7.95 22.05 10.50 ;
        RECT  21.25 4.05 22.15 4.95 ;
        RECT  21.25 7.95 22.15 8.90 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  24.05 2.70 24.75 4.50 ;
        RECT  24.25 2.70 24.75 10.50 ;
        RECT  24.05 7.95 24.75 10.50 ;
        RECT  24.05 7.95 24.95 8.95 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  40.85 5.40 41.75 6.30 ;
        RECT  40.30 5.60 41.75 6.30 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  42.25 5.40 43.15 6.30 ;
        END
    END J
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.25 6.65 2.55 7.35 ;
        RECT  1.65 6.65 2.55 7.65 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.30 2.50 11.00 ;
        RECT  4.05 7.95 4.75 11.00 ;
        RECT  9.80 8.10 10.50 11.00 ;
        RECT  12.30 9.55 13.00 11.00 ;
        RECT  17.15 9.05 17.85 11.00 ;
        RECT  19.85 9.15 20.55 11.00 ;
        RECT  22.70 7.65 23.40 11.00 ;
        RECT  27.20 7.10 27.90 11.00 ;
        RECT  39.40 7.80 40.10 11.00 ;
        RECT  42.25 7.10 42.95 11.00 ;
        RECT  0.00 11.00 44.80 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.90 2.00 1.70 3.20 ;
        RECT  4.05 2.00 4.75 4.85 ;
        RECT  8.50 2.00 9.00 4.25 ;
        RECT  9.90 3.75 10.60 4.95 ;
        RECT  8.50 3.75 13.60 4.25 ;
        RECT  12.90 3.75 13.60 5.00 ;
        RECT  17.60 4.25 18.30 5.00 ;
        RECT  18.45 2.00 18.95 4.75 ;
        RECT  17.60 4.25 18.95 4.75 ;
        RECT  22.70 2.00 23.40 4.50 ;
        RECT  27.20 2.00 27.90 4.45 ;
        RECT  34.20 2.00 34.90 4.15 ;
        RECT  42.25 2.00 42.95 4.45 ;
        RECT  0.00 0.00 44.80 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.25 5.35 0.75 10.25 ;
        RECT  0.25 9.55 1.15 10.25 ;
        RECT  1.00 3.80 1.80 5.85 ;
        RECT  0.25 5.35 1.80 5.85 ;
        RECT  2.70 4.20 3.55 4.90 ;
        RECT  3.05 4.20 3.55 8.85 ;
        RECT  2.70 8.15 3.55 8.85 ;
        RECT  3.05 5.55 6.35 6.05 ;
        RECT  5.35 3.20 5.85 6.05 ;
        RECT  5.85 5.55 6.35 7.40 ;
        RECT  5.85 6.70 6.55 7.40 ;
        RECT  6.40 4.20 7.55 4.90 ;
        RECT  6.85 3.00 7.55 3.70 ;
        RECT  5.35 3.20 7.55 3.70 ;
        RECT  7.05 4.20 7.55 9.25 ;
        RECT  6.40 8.55 8.00 9.25 ;
        RECT  9.35 5.65 10.05 6.35 ;
        RECT  10.35 6.90 11.05 7.60 ;
        RECT  7.05 7.10 11.05 7.60 ;
        RECT  11.40 4.75 12.10 6.15 ;
        RECT  9.35 5.65 12.10 6.15 ;
        RECT  11.60 4.75 12.10 8.85 ;
        RECT  11.15 8.10 12.10 8.85 ;
        RECT  15.25 4.30 15.50 9.85 ;
        RECT  14.80 7.15 15.50 9.85 ;
        RECT  15.25 4.30 15.75 7.65 ;
        RECT  15.25 4.30 15.95 5.00 ;
        RECT  16.95 5.95 17.65 6.70 ;
        RECT  18.50 8.15 19.20 9.85 ;
        RECT  19.00 6.95 19.70 7.65 ;
        RECT  14.80 7.15 19.70 7.65 ;
        RECT  20.20 4.35 20.65 8.65 ;
        RECT  19.95 4.35 20.65 6.45 ;
        RECT  20.20 5.95 20.70 8.65 ;
        RECT  18.50 8.15 20.70 8.65 ;
        RECT  23.05 5.75 23.75 6.45 ;
        RECT  16.95 5.95 23.75 6.45 ;
        RECT  25.50 2.55 26.35 3.25 ;
        RECT  25.80 2.55 26.35 8.90 ;
        RECT  25.80 3.75 26.55 4.45 ;
        RECT  25.80 7.10 26.60 8.90 ;
        RECT  28.55 3.75 29.25 4.45 ;
        RECT  28.55 7.10 29.25 8.90 ;
        RECT  28.55 3.95 30.15 4.45 ;
        RECT  29.65 3.95 30.15 7.60 ;
        RECT  28.55 7.10 30.15 7.60 ;
        RECT  30.20 9.75 30.90 10.45 ;
        RECT  30.65 4.60 31.35 5.30 ;
        RECT  31.50 6.80 32.00 9.45 ;
        RECT  31.30 7.75 32.00 9.45 ;
        RECT  31.65 3.70 32.35 5.10 ;
        RECT  32.65 7.80 33.35 10.45 ;
        RECT  30.20 9.95 33.35 10.45 ;
        RECT  34.00 6.80 34.70 10.45 ;
        RECT  35.35 7.80 36.05 10.45 ;
        RECT  31.50 6.80 37.20 7.30 ;
        RECT  36.70 6.80 37.20 9.45 ;
        RECT  36.70 7.75 37.40 9.45 ;
        RECT  37.40 5.60 38.10 6.30 ;
        RECT  29.65 5.80 38.10 6.30 ;
        RECT  37.70 3.45 38.20 5.10 ;
        RECT  30.65 4.60 38.20 5.10 ;
        RECT  38.05 7.80 38.75 10.45 ;
        RECT  38.25 6.80 38.75 10.45 ;
        RECT  35.35 9.95 38.75 10.45 ;
        RECT  37.70 3.45 39.30 4.15 ;
        RECT  38.25 6.80 41.25 7.30 ;
        RECT  40.75 6.80 41.25 10.50 ;
        RECT  40.75 7.80 41.45 10.50 ;
        RECT  43.65 3.75 44.15 10.50 ;
        RECT  43.65 3.75 44.35 4.45 ;
        RECT  43.65 7.10 44.35 10.50 ;
        RECT  43.65 9.80 44.50 10.50 ;
        LAYER V1M ;
        RECT  21.20 7.95 22.20 8.95 ;
        RECT  21.20 4.05 22.20 5.05 ;
    END
END SJKRRX2
MACRO SJKRRX4
    CLASS CORE ;
    FOREIGN SJKRRX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 47.60 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  31.05 5.40 31.95 6.30 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  29.65 5.40 30.55 6.30 ;
        END
    END SD
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  9.50 2.55 10.20 3.25 ;
        RECT  15.65 2.70 16.55 3.70 ;
        RECT  17.15 2.55 17.85 3.25 ;
        RECT  9.50 2.70 17.85 3.25 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M2M ;
        RECT  22.80 4.10 23.40 9.00 ;
        RECT  22.70 4.10 23.50 4.90 ;
        RECT  22.70 7.90 23.50 9.00 ;
        LAYER M1M ;
        RECT  22.80 2.75 23.50 4.95 ;
        RECT  22.80 7.95 23.50 10.50 ;
        RECT  22.65 4.05 23.55 4.95 ;
        RECT  22.65 7.95 23.55 8.90 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  25.50 2.70 26.20 4.50 ;
        RECT  25.70 2.70 26.20 10.50 ;
        RECT  25.50 7.95 26.20 10.50 ;
        RECT  25.45 7.95 26.35 8.95 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  43.65 5.40 44.55 6.30 ;
        RECT  43.10 5.60 44.55 6.30 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  45.05 5.40 45.95 6.30 ;
        END
    END J
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.25 6.65 2.55 7.35 ;
        RECT  1.65 6.65 2.55 7.65 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.30 2.50 11.00 ;
        RECT  4.05 7.95 4.75 11.00 ;
        RECT  9.80 8.10 10.50 11.00 ;
        RECT  12.30 9.55 13.00 11.00 ;
        RECT  17.15 9.05 17.85 11.00 ;
        RECT  19.85 9.15 20.55 11.00 ;
        RECT  21.45 7.65 22.15 11.00 ;
        RECT  24.15 7.65 24.85 11.00 ;
        RECT  26.85 7.65 27.55 11.00 ;
        RECT  30.00 7.10 30.70 11.00 ;
        RECT  42.20 7.80 42.90 11.00 ;
        RECT  45.05 7.10 45.75 11.00 ;
        RECT  0.00 11.00 47.60 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.90 2.00 1.70 3.20 ;
        RECT  4.05 2.00 4.75 4.85 ;
        RECT  8.50 2.00 9.00 4.25 ;
        RECT  9.90 3.75 10.60 4.95 ;
        RECT  8.50 3.75 13.60 4.25 ;
        RECT  12.90 3.75 13.60 5.00 ;
        RECT  17.60 4.25 18.30 5.00 ;
        RECT  18.45 2.00 18.95 4.75 ;
        RECT  17.60 4.25 18.95 4.75 ;
        RECT  21.45 2.00 22.15 4.50 ;
        RECT  24.15 2.00 24.85 4.50 ;
        RECT  26.85 2.00 27.55 4.50 ;
        RECT  30.00 2.00 30.70 4.45 ;
        RECT  37.00 2.00 37.70 4.15 ;
        RECT  45.05 2.00 45.75 4.45 ;
        RECT  0.00 0.00 47.60 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.25 5.35 0.75 10.25 ;
        RECT  0.25 9.55 1.15 10.25 ;
        RECT  1.00 3.80 1.80 5.85 ;
        RECT  0.25 5.35 1.80 5.85 ;
        RECT  2.70 4.20 3.55 4.90 ;
        RECT  3.05 4.20 3.55 8.85 ;
        RECT  2.70 8.15 3.55 8.85 ;
        RECT  3.05 5.55 6.35 6.05 ;
        RECT  5.35 3.20 5.85 6.05 ;
        RECT  5.85 5.55 6.35 7.40 ;
        RECT  5.85 6.70 6.55 7.40 ;
        RECT  6.40 4.20 7.55 4.90 ;
        RECT  6.85 3.00 7.55 3.70 ;
        RECT  5.35 3.20 7.55 3.70 ;
        RECT  7.05 4.20 7.55 9.25 ;
        RECT  6.40 8.55 8.00 9.25 ;
        RECT  9.35 5.65 10.05 6.35 ;
        RECT  10.35 6.90 11.05 7.60 ;
        RECT  7.05 7.10 11.05 7.60 ;
        RECT  11.40 4.75 12.10 6.15 ;
        RECT  9.35 5.65 12.10 6.15 ;
        RECT  11.60 4.75 12.10 8.85 ;
        RECT  11.15 8.10 12.10 8.85 ;
        RECT  15.25 4.30 15.50 9.85 ;
        RECT  14.80 7.15 15.50 9.85 ;
        RECT  15.25 4.30 15.75 7.65 ;
        RECT  15.25 4.30 15.95 5.00 ;
        RECT  16.95 5.95 17.65 6.70 ;
        RECT  18.50 8.15 19.20 9.85 ;
        RECT  19.00 6.95 19.70 7.65 ;
        RECT  14.80 7.15 19.70 7.65 ;
        RECT  20.20 4.35 20.65 8.65 ;
        RECT  19.95 4.35 20.65 6.45 ;
        RECT  20.20 5.95 20.70 8.65 ;
        RECT  18.50 8.15 20.70 8.65 ;
        RECT  24.50 5.75 25.20 6.45 ;
        RECT  16.95 5.95 25.20 6.45 ;
        RECT  28.30 2.55 29.15 3.25 ;
        RECT  28.60 2.55 29.15 8.90 ;
        RECT  28.60 3.75 29.35 4.45 ;
        RECT  28.60 7.10 29.40 8.90 ;
        RECT  31.35 3.75 32.05 4.45 ;
        RECT  31.35 7.10 32.05 8.90 ;
        RECT  31.35 3.95 32.95 4.45 ;
        RECT  32.45 3.95 32.95 7.60 ;
        RECT  31.35 7.10 32.95 7.60 ;
        RECT  33.00 9.75 33.70 10.45 ;
        RECT  33.45 4.60 34.15 5.30 ;
        RECT  34.30 6.80 34.80 9.45 ;
        RECT  34.10 7.75 34.80 9.45 ;
        RECT  34.45 3.70 35.15 5.10 ;
        RECT  35.45 7.80 36.15 10.45 ;
        RECT  33.00 9.95 36.15 10.45 ;
        RECT  36.80 6.80 37.50 10.45 ;
        RECT  38.15 7.80 38.85 10.45 ;
        RECT  34.30 6.80 40.00 7.30 ;
        RECT  39.50 6.80 40.00 9.45 ;
        RECT  39.50 7.75 40.20 9.45 ;
        RECT  40.20 5.60 40.90 6.30 ;
        RECT  32.45 5.80 40.90 6.30 ;
        RECT  40.50 3.45 41.00 5.10 ;
        RECT  33.45 4.60 41.00 5.10 ;
        RECT  40.85 7.80 41.55 10.45 ;
        RECT  41.05 6.80 41.55 10.45 ;
        RECT  38.15 9.95 41.55 10.45 ;
        RECT  40.50 3.45 42.10 4.15 ;
        RECT  41.05 6.80 44.05 7.30 ;
        RECT  43.55 6.80 44.05 10.50 ;
        RECT  43.55 7.80 44.25 10.50 ;
        RECT  46.45 3.75 46.95 10.50 ;
        RECT  46.45 3.75 47.15 4.45 ;
        RECT  46.45 7.10 47.15 10.50 ;
        RECT  46.45 9.80 47.30 10.50 ;
        LAYER V1M ;
        RECT  22.60 7.95 23.60 8.95 ;
        RECT  22.60 4.05 23.60 5.05 ;
    END
END SJKRRX4
MACRO SJKRSX1
    CLASS CORE ;
    FOREIGN SJKRSX1 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 43.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  11.45 7.05 12.15 7.75 ;
        RECT  12.85 6.70 13.75 7.60 ;
        RECT  13.25 5.45 13.75 7.60 ;
        RECT  11.45 7.05 13.75 7.60 ;
        RECT  13.90 5.25 14.60 5.95 ;
        RECT  13.25 5.45 14.60 5.95 ;
        END
    END SN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  26.85 5.40 27.75 6.30 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  25.45 5.40 26.35 6.30 ;
        END
    END SD
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M2M ;
        RECT  20.00 4.35 20.60 7.70 ;
        RECT  19.90 4.35 20.70 5.15 ;
        RECT  19.90 6.60 20.70 7.70 ;
        LAYER M1M ;
        RECT  19.85 6.70 20.75 7.60 ;
        RECT  20.05 3.75 20.75 5.20 ;
        RECT  19.85 4.30 20.75 5.20 ;
        RECT  20.05 6.70 20.75 8.90 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  22.75 3.75 23.45 4.45 ;
        RECT  22.95 3.75 23.45 8.90 ;
        RECT  22.75 6.70 23.45 8.90 ;
        RECT  22.65 6.70 23.55 7.60 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  39.45 5.40 40.35 6.30 ;
        RECT  38.90 5.60 40.35 6.30 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  40.85 5.40 41.75 6.30 ;
        END
    END J
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.25 6.65 2.55 7.35 ;
        RECT  1.65 6.65 2.55 7.65 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.30 2.50 11.00 ;
        RECT  4.05 7.95 4.75 11.00 ;
        RECT  8.75 7.90 9.45 11.00 ;
        RECT  8.00 10.45 9.60 11.00 ;
        RECT  12.05 8.70 12.75 11.00 ;
        RECT  17.05 7.10 17.75 11.00 ;
        RECT  21.40 7.10 22.10 11.00 ;
        RECT  19.50 10.45 23.50 11.00 ;
        RECT  25.80 7.10 26.50 11.00 ;
        RECT  38.00 7.80 38.70 11.00 ;
        RECT  40.85 7.10 41.55 11.00 ;
        RECT  0.00 11.00 43.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.90 2.00 1.70 3.20 ;
        RECT  4.05 2.00 4.75 4.85 ;
        RECT  8.15 2.00 9.75 3.15 ;
        RECT  9.05 2.00 9.75 4.90 ;
        RECT  11.20 2.00 11.90 3.25 ;
        RECT  17.05 2.00 17.75 3.95 ;
        RECT  21.40 2.00 22.10 4.40 ;
        RECT  25.80 2.00 26.50 4.45 ;
        RECT  32.80 2.00 33.50 4.15 ;
        RECT  40.85 2.00 41.55 4.45 ;
        RECT  0.00 0.00 43.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.25 5.35 0.75 10.25 ;
        RECT  0.25 9.55 1.20 10.25 ;
        RECT  1.00 3.80 1.80 5.85 ;
        RECT  0.25 5.35 1.80 5.85 ;
        RECT  2.70 4.20 3.55 4.90 ;
        RECT  3.05 4.20 3.55 8.85 ;
        RECT  2.70 8.15 3.55 8.85 ;
        RECT  3.05 5.55 6.35 6.05 ;
        RECT  5.35 3.20 5.85 6.05 ;
        RECT  5.85 5.55 6.35 7.40 ;
        RECT  5.85 6.70 6.55 7.40 ;
        RECT  6.40 4.20 7.10 4.90 ;
        RECT  6.40 4.40 7.55 4.90 ;
        RECT  7.05 4.20 7.10 9.55 ;
        RECT  6.40 7.90 7.10 9.55 ;
        RECT  6.85 3.00 7.55 3.70 ;
        RECT  5.35 3.20 7.55 3.70 ;
        RECT  7.05 4.40 7.55 8.40 ;
        RECT  6.40 7.90 7.55 8.40 ;
        RECT  8.30 5.45 9.00 6.15 ;
        RECT  7.05 6.70 9.95 7.20 ;
        RECT  9.25 6.70 9.95 7.40 ;
        RECT  8.30 5.45 10.95 5.95 ;
        RECT  10.45 4.35 10.95 9.45 ;
        RECT  10.45 8.75 11.25 9.45 ;
        RECT  11.55 4.15 12.25 4.85 ;
        RECT  10.45 4.35 12.25 4.85 ;
        RECT  13.70 3.30 14.40 4.00 ;
        RECT  13.70 3.45 15.60 4.00 ;
        RECT  14.55 7.20 15.10 10.50 ;
        RECT  14.40 8.70 15.10 10.50 ;
        RECT  15.10 3.45 15.60 7.90 ;
        RECT  14.55 7.20 15.60 7.90 ;
        RECT  16.60 4.45 17.30 5.15 ;
        RECT  17.40 5.70 18.10 6.40 ;
        RECT  15.10 5.90 18.10 6.40 ;
        RECT  18.40 3.25 19.10 3.95 ;
        RECT  16.60 4.45 19.10 4.95 ;
        RECT  18.55 7.10 19.25 8.90 ;
        RECT  18.75 3.25 19.10 9.95 ;
        RECT  18.60 3.25 19.10 8.90 ;
        RECT  18.75 7.10 19.25 9.95 ;
        RECT  18.75 9.25 19.60 9.95 ;
        RECT  21.75 5.50 22.45 6.20 ;
        RECT  18.60 5.70 22.45 6.20 ;
        RECT  24.10 2.55 24.95 3.25 ;
        RECT  24.40 2.55 24.95 8.90 ;
        RECT  24.40 3.75 25.15 4.45 ;
        RECT  24.40 7.10 25.20 8.90 ;
        RECT  27.15 3.75 27.85 4.45 ;
        RECT  27.15 7.10 27.85 8.90 ;
        RECT  27.15 3.95 28.75 4.45 ;
        RECT  28.25 3.95 28.75 7.60 ;
        RECT  27.15 7.10 28.75 7.60 ;
        RECT  28.80 9.75 29.50 10.45 ;
        RECT  29.25 4.60 29.95 5.30 ;
        RECT  30.10 6.80 30.60 9.45 ;
        RECT  29.90 7.75 30.60 9.45 ;
        RECT  30.25 3.70 30.95 5.10 ;
        RECT  31.25 7.80 31.95 10.45 ;
        RECT  28.80 9.95 31.95 10.45 ;
        RECT  32.60 6.80 33.30 10.45 ;
        RECT  33.95 7.80 34.65 10.45 ;
        RECT  30.10 6.80 35.80 7.30 ;
        RECT  35.30 6.80 35.80 9.45 ;
        RECT  35.30 7.75 36.00 9.45 ;
        RECT  36.00 5.60 36.70 6.30 ;
        RECT  28.25 5.80 36.70 6.30 ;
        RECT  36.30 3.45 36.80 5.10 ;
        RECT  29.25 4.60 36.80 5.10 ;
        RECT  36.65 7.80 37.35 10.45 ;
        RECT  36.85 6.80 37.35 10.45 ;
        RECT  33.95 9.95 37.35 10.45 ;
        RECT  36.30 3.45 37.90 4.15 ;
        RECT  36.85 6.80 39.85 7.30 ;
        RECT  39.35 6.80 39.85 10.50 ;
        RECT  39.35 7.80 40.05 10.50 ;
        RECT  42.25 3.75 42.75 10.50 ;
        RECT  42.25 3.75 42.95 4.45 ;
        RECT  42.25 7.10 42.95 10.50 ;
        RECT  42.25 9.80 43.10 10.50 ;
        LAYER V1M ;
        RECT  19.80 6.65 20.80 7.65 ;
        RECT  19.80 4.05 20.80 5.05 ;
    END
END SJKRSX1
MACRO SJKRSX2
    CLASS CORE ;
    FOREIGN SJKRSX2 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 43.40 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  11.45 7.05 12.15 7.75 ;
        RECT  12.85 6.70 13.75 7.60 ;
        RECT  13.25 5.45 13.75 7.60 ;
        RECT  11.45 7.05 13.75 7.60 ;
        RECT  13.90 5.25 14.60 5.95 ;
        RECT  13.25 5.45 14.60 5.95 ;
        END
    END SN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  26.85 5.40 27.75 6.30 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  25.45 5.40 26.35 6.30 ;
        END
    END SD
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M2M ;
        RECT  20.00 4.35 20.60 7.70 ;
        RECT  19.90 4.35 20.70 5.15 ;
        RECT  19.90 6.60 20.70 7.70 ;
        LAYER M1M ;
        RECT  19.85 6.70 20.75 7.60 ;
        RECT  20.05 2.70 20.75 5.20 ;
        RECT  19.85 4.30 20.75 5.20 ;
        RECT  20.05 6.70 20.75 10.50 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  22.75 2.70 23.45 4.50 ;
        RECT  22.95 2.70 23.45 10.50 ;
        RECT  22.75 6.70 23.45 10.50 ;
        RECT  22.65 6.70 23.55 7.60 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  39.45 5.40 40.35 6.30 ;
        RECT  38.90 5.60 40.35 6.30 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  40.85 5.40 41.75 6.30 ;
        END
    END J
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.25 6.65 2.55 7.35 ;
        RECT  1.65 6.65 2.55 7.65 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.30 2.50 11.00 ;
        RECT  4.05 7.95 4.75 11.00 ;
        RECT  8.75 7.90 9.45 11.00 ;
        RECT  8.00 10.45 9.60 11.00 ;
        RECT  12.05 8.70 12.75 11.00 ;
        RECT  17.05 7.10 17.75 11.00 ;
        RECT  21.40 7.10 22.10 11.00 ;
        RECT  25.80 7.10 26.50 11.00 ;
        RECT  38.00 7.80 38.70 11.00 ;
        RECT  40.85 7.10 41.55 11.00 ;
        RECT  0.00 11.00 43.40 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.90 2.00 1.70 3.20 ;
        RECT  4.05 2.00 4.75 4.85 ;
        RECT  8.15 2.00 9.75 3.15 ;
        RECT  9.05 2.00 9.75 4.90 ;
        RECT  11.20 2.00 11.90 3.25 ;
        RECT  17.05 2.00 17.75 3.95 ;
        RECT  21.40 2.00 22.10 4.50 ;
        RECT  25.80 2.00 26.50 4.45 ;
        RECT  32.80 2.00 33.50 4.15 ;
        RECT  40.85 2.00 41.55 4.45 ;
        RECT  0.00 0.00 43.40 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.25 5.35 0.75 10.25 ;
        RECT  0.25 9.55 1.20 10.25 ;
        RECT  1.00 3.80 1.80 5.85 ;
        RECT  0.25 5.35 1.80 5.85 ;
        RECT  2.70 4.20 3.55 4.90 ;
        RECT  3.05 4.20 3.55 8.85 ;
        RECT  2.70 8.15 3.55 8.85 ;
        RECT  3.05 5.55 6.35 6.05 ;
        RECT  5.35 3.20 5.85 6.05 ;
        RECT  5.85 5.55 6.35 7.40 ;
        RECT  5.85 6.70 6.55 7.40 ;
        RECT  6.40 4.20 7.10 4.90 ;
        RECT  6.40 4.40 7.55 4.90 ;
        RECT  7.05 4.20 7.10 9.55 ;
        RECT  6.40 7.90 7.10 9.55 ;
        RECT  6.85 3.00 7.55 3.70 ;
        RECT  5.35 3.20 7.55 3.70 ;
        RECT  7.05 4.40 7.55 8.40 ;
        RECT  6.40 7.90 7.55 8.40 ;
        RECT  8.30 5.45 9.00 6.15 ;
        RECT  7.05 6.70 9.95 7.20 ;
        RECT  9.25 6.70 9.95 7.40 ;
        RECT  8.30 5.45 10.95 5.95 ;
        RECT  10.45 4.35 10.95 9.45 ;
        RECT  10.45 8.75 11.25 9.45 ;
        RECT  11.55 4.15 12.25 4.85 ;
        RECT  10.45 4.35 12.25 4.85 ;
        RECT  13.70 3.30 14.40 4.00 ;
        RECT  13.70 3.45 15.60 4.00 ;
        RECT  14.55 7.20 15.10 10.50 ;
        RECT  14.40 8.70 15.10 10.50 ;
        RECT  15.10 3.45 15.60 7.90 ;
        RECT  14.55 7.20 15.60 7.90 ;
        RECT  16.60 4.45 17.30 5.15 ;
        RECT  17.40 5.70 18.10 6.40 ;
        RECT  15.10 5.90 18.10 6.40 ;
        RECT  18.40 3.25 19.10 3.95 ;
        RECT  16.60 4.45 19.10 4.95 ;
        RECT  18.55 7.10 19.25 8.90 ;
        RECT  18.75 3.25 19.10 10.50 ;
        RECT  18.60 3.25 19.10 8.90 ;
        RECT  18.75 7.10 19.25 10.50 ;
        RECT  18.75 9.80 19.55 10.50 ;
        RECT  21.75 5.50 22.45 6.20 ;
        RECT  18.60 5.70 22.45 6.20 ;
        RECT  24.10 2.55 24.95 3.25 ;
        RECT  24.40 2.55 24.95 8.90 ;
        RECT  24.40 3.75 25.15 4.45 ;
        RECT  24.40 7.10 25.20 8.90 ;
        RECT  27.15 3.75 27.85 4.45 ;
        RECT  27.15 7.10 27.85 8.90 ;
        RECT  27.15 3.95 28.75 4.45 ;
        RECT  28.25 3.95 28.75 7.60 ;
        RECT  27.15 7.10 28.75 7.60 ;
        RECT  28.80 9.75 29.50 10.45 ;
        RECT  29.25 4.60 29.95 5.30 ;
        RECT  30.10 6.80 30.60 9.45 ;
        RECT  29.90 7.75 30.60 9.45 ;
        RECT  30.25 3.70 30.95 5.10 ;
        RECT  31.25 7.80 31.95 10.45 ;
        RECT  28.80 9.95 31.95 10.45 ;
        RECT  32.60 6.80 33.30 10.45 ;
        RECT  33.95 7.80 34.65 10.45 ;
        RECT  30.10 6.80 35.80 7.30 ;
        RECT  35.30 6.80 35.80 9.45 ;
        RECT  35.30 7.75 36.00 9.45 ;
        RECT  36.00 5.60 36.70 6.30 ;
        RECT  28.25 5.80 36.70 6.30 ;
        RECT  36.30 3.45 36.80 5.10 ;
        RECT  29.25 4.60 36.80 5.10 ;
        RECT  36.65 7.80 37.35 10.45 ;
        RECT  36.85 6.80 37.35 10.45 ;
        RECT  33.95 9.95 37.35 10.45 ;
        RECT  36.30 3.45 37.90 4.15 ;
        RECT  36.85 6.80 39.85 7.30 ;
        RECT  39.35 6.80 39.85 10.50 ;
        RECT  39.35 7.80 40.05 10.50 ;
        RECT  42.25 3.75 42.75 10.50 ;
        RECT  42.25 3.75 42.95 4.45 ;
        RECT  42.25 7.10 42.95 10.50 ;
        RECT  42.25 9.80 43.10 10.50 ;
        LAYER V1M ;
        RECT  19.80 6.65 20.80 7.65 ;
        RECT  19.80 4.05 20.80 5.05 ;
    END
END SJKRSX2
MACRO SJKRSX4
    CLASS CORE ;
    FOREIGN SJKRSX4 0.00 0.00  ;
    ORIGIN 0.00 0.00 ;
    SIZE 46.20 BY 13.00 ;
    SYMMETRY x y r90 ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.40 ;
        PORT
        LAYER M1M ;
        RECT  11.45 7.05 12.15 7.75 ;
        RECT  12.85 6.70 13.75 7.60 ;
        RECT  13.25 5.45 13.75 7.60 ;
        RECT  11.45 7.05 13.75 7.60 ;
        RECT  13.90 5.25 14.60 5.95 ;
        RECT  13.25 5.45 14.60 5.95 ;
        END
    END SN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.45 ;
        PORT
        LAYER M1M ;
        RECT  29.65 5.40 30.55 6.30 ;
        END
    END SE
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  28.25 5.40 29.15 6.30 ;
        END
    END SD
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M2M ;
        RECT  21.40 4.10 22.00 9.00 ;
        RECT  21.30 4.10 22.10 4.90 ;
        RECT  21.30 7.90 22.10 9.00 ;
        LAYER M1M ;
        RECT  21.40 2.75 22.10 4.95 ;
        RECT  21.40 7.95 22.10 10.50 ;
        RECT  21.25 4.05 22.15 4.95 ;
        RECT  21.25 7.95 22.15 8.90 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.0 ;
        PORT
        LAYER M1M ;
        RECT  24.10 2.70 24.80 4.50 ;
        RECT  24.30 2.70 24.80 10.50 ;
        RECT  24.10 7.95 24.80 10.50 ;
        RECT  24.05 7.95 24.95 8.95 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.57 ;
        PORT
        LAYER M1M ;
        RECT  42.25 5.40 43.15 6.30 ;
        RECT  41.70 5.60 43.15 6.30 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  43.65 5.40 44.55 6.30 ;
        END
    END J
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.05 ;
        PORT
        LAYER M1M ;
        RECT  1.25 6.65 2.55 7.35 ;
        RECT  1.65 6.65 2.55 7.65 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  1.80 10.30 2.50 11.00 ;
        RECT  4.05 7.95 4.75 11.00 ;
        RECT  8.75 7.90 9.45 11.00 ;
        RECT  8.00 10.45 9.60 11.00 ;
        RECT  12.05 8.70 12.75 11.00 ;
        RECT  17.05 7.10 17.75 11.00 ;
        RECT  20.05 7.65 20.75 11.00 ;
        RECT  22.75 7.65 23.45 11.00 ;
        RECT  25.45 7.65 26.15 11.00 ;
        RECT  28.60 7.10 29.30 11.00 ;
        RECT  40.80 7.80 41.50 11.00 ;
        RECT  43.65 7.10 44.35 11.00 ;
        RECT  0.00 11.00 46.20 13.00 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1M ;
        RECT  0.90 2.00 1.70 3.20 ;
        RECT  4.05 2.00 4.75 4.85 ;
        RECT  8.15 2.00 9.75 3.15 ;
        RECT  9.05 2.00 9.75 4.90 ;
        RECT  11.20 2.00 11.90 3.25 ;
        RECT  17.05 2.00 17.75 3.95 ;
        RECT  20.05 2.00 20.75 4.50 ;
        RECT  22.75 2.00 23.45 4.50 ;
        RECT  25.45 2.00 26.15 4.50 ;
        RECT  28.60 2.00 29.30 4.45 ;
        RECT  35.60 2.00 36.30 4.15 ;
        RECT  43.65 2.00 44.35 4.45 ;
        RECT  0.00 0.00 46.20 2.00 ;
        END
    END gnd!
    OBS
        LAYER M1M ;
        RECT  0.25 5.35 0.75 10.25 ;
        RECT  0.25 9.55 1.20 10.25 ;
        RECT  1.00 3.80 1.80 5.85 ;
        RECT  0.25 5.35 1.80 5.85 ;
        RECT  2.70 4.20 3.55 4.90 ;
        RECT  3.05 4.20 3.55 8.85 ;
        RECT  2.70 8.15 3.55 8.85 ;
        RECT  3.05 5.55 6.35 6.05 ;
        RECT  5.35 3.20 5.85 6.05 ;
        RECT  5.85 5.55 6.35 7.40 ;
        RECT  5.85 6.70 6.55 7.40 ;
        RECT  6.40 4.20 7.10 4.90 ;
        RECT  6.40 4.40 7.55 4.90 ;
        RECT  7.05 4.20 7.10 9.55 ;
        RECT  6.40 7.90 7.10 9.55 ;
        RECT  6.85 3.00 7.55 3.70 ;
        RECT  5.35 3.20 7.55 3.70 ;
        RECT  7.05 4.40 7.55 8.40 ;
        RECT  6.40 7.90 7.55 8.40 ;
        RECT  8.30 5.45 9.00 6.15 ;
        RECT  7.05 6.70 9.95 7.20 ;
        RECT  9.25 6.70 9.95 7.40 ;
        RECT  8.30 5.45 10.95 5.95 ;
        RECT  10.45 4.35 10.95 9.45 ;
        RECT  10.45 8.75 11.25 9.45 ;
        RECT  11.55 4.15 12.25 4.85 ;
        RECT  10.45 4.35 12.25 4.85 ;
        RECT  13.70 3.30 14.40 4.00 ;
        RECT  13.70 3.45 15.60 4.00 ;
        RECT  14.55 7.20 15.10 10.50 ;
        RECT  14.40 8.70 15.10 10.50 ;
        RECT  15.10 3.45 15.60 7.90 ;
        RECT  14.55 7.20 15.60 7.90 ;
        RECT  16.60 4.45 17.30 5.15 ;
        RECT  17.40 5.70 18.10 6.40 ;
        RECT  15.10 5.90 18.10 6.40 ;
        RECT  18.40 3.25 19.10 3.95 ;
        RECT  16.60 4.45 19.10 4.95 ;
        RECT  18.55 7.10 19.25 8.90 ;
        RECT  18.75 3.25 19.10 10.50 ;
        RECT  18.60 3.25 19.10 8.90 ;
        RECT  18.75 7.10 19.25 10.50 ;
        RECT  18.75 9.80 19.55 10.50 ;
        RECT  23.10 5.75 23.80 6.45 ;
        RECT  18.60 5.95 23.80 6.45 ;
        RECT  26.90 2.55 27.75 3.25 ;
        RECT  27.20 2.55 27.75 8.90 ;
        RECT  27.20 3.75 27.95 4.45 ;
        RECT  27.20 7.10 28.00 8.90 ;
        RECT  29.95 3.75 30.65 4.45 ;
        RECT  29.95 7.10 30.65 8.90 ;
        RECT  29.95 3.95 31.55 4.45 ;
        RECT  31.05 3.95 31.55 7.60 ;
        RECT  29.95 7.10 31.55 7.60 ;
        RECT  31.60 9.75 32.30 10.45 ;
        RECT  32.05 4.60 32.75 5.30 ;
        RECT  32.90 6.80 33.40 9.45 ;
        RECT  32.70 7.75 33.40 9.45 ;
        RECT  33.05 3.70 33.75 5.10 ;
        RECT  34.05 7.80 34.75 10.45 ;
        RECT  31.60 9.95 34.75 10.45 ;
        RECT  35.40 6.80 36.10 10.45 ;
        RECT  36.75 7.80 37.45 10.45 ;
        RECT  32.90 6.80 38.60 7.30 ;
        RECT  38.10 6.80 38.60 9.45 ;
        RECT  38.10 7.75 38.80 9.45 ;
        RECT  38.80 5.60 39.50 6.30 ;
        RECT  31.05 5.80 39.50 6.30 ;
        RECT  39.10 3.45 39.60 5.10 ;
        RECT  32.05 4.60 39.60 5.10 ;
        RECT  39.45 7.80 40.15 10.45 ;
        RECT  39.65 6.80 40.15 10.45 ;
        RECT  36.75 9.95 40.15 10.45 ;
        RECT  39.10 3.45 40.70 4.15 ;
        RECT  39.65 6.80 42.65 7.30 ;
        RECT  42.15 6.80 42.65 10.50 ;
        RECT  42.15 7.80 42.85 10.50 ;
        RECT  45.05 3.75 45.55 10.50 ;
        RECT  45.05 3.75 45.75 4.45 ;
        RECT  45.05 7.10 45.75 10.50 ;
        RECT  45.05 9.80 45.90 10.50 ;
        LAYER V1M ;
        RECT  21.20 7.95 22.20 8.95 ;
        RECT  21.20 4.05 22.20 5.05 ;
    END
END SJKRSX4
END LIBRARY
